* SPICE3 file created from TWOBIT_FLASH_ADC_0.ext - technology: sky130A
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.subckt TWOBIT_FLASH_ADC GND VCC C3 C2 C1 VREF2 VREF3 VREF1 BIAS INP
X0 GND COMP_PG0_2_0_1680520037_0/m1_2720_1484# C1 GND sky130_fd_pr__nfet_01v8 ad=8.1648e+12p pd=7.992e+07u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X1 C1 COMP_PG0_2_0_1680520037_0/m1_2720_1484# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 GND COMP_PG0_2_0_1680520037_0/m1_2720_1484# C1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 C1 COMP_PG0_2_0_1680520037_0/m1_2720_1484# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 C1 COMP_PG0_2_0_1680520037_0/m1_2720_1484# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=9.576e+12p ps=9.336e+07u w=840000u l=150000u
X5 VCC COMP_PG0_2_0_1680520037_0/m1_2720_1484# C1 VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 C1 COMP_PG0_2_0_1680520037_0/m1_2720_1484# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 VCC COMP_PG0_2_0_1680520037_0/m1_2720_1484# C1 VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 GND COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_2720_1484# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X9 COMP_PG0_2_0_1680520037_0/m1_2720_1484# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 GND COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_2720_1484# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 COMP_PG0_2_0_1680520037_0/m1_2720_1484# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 GND COMP_PG0_2_0_1680520037_0/m1_1172_1316# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X13 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_1172_1316# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 GND COMP_PG0_2_0_1680520037_0/m1_1172_1316# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_1172_1316# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 COMP_PG0_2_0_1680520037_0/m1_2720_1484# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X17 VCC COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_2720_1484# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18 COMP_PG0_2_0_1680520037_0/m1_2720_1484# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 VCC COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_2720_1484# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_1172_1316# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X21 VCC COMP_PG0_2_0_1680520037_0/m1_1172_1316# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_1172_1316# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 VCC COMP_PG0_2_0_1680520037_0/m1_1172_1316# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24 COMP_PG0_2_0_1680520037_0/m1_688_1652# INP COMP_PG0_2_0_1680520037_0/m1_1172_1316# GND sky130_fd_pr__nfet_01v8 ad=1.8312e+12p pd=1.78e+07u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X25 COMP_PG0_2_0_1680520037_0/m1_1172_1316# INP COMP_PG0_2_0_1680520037_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 COMP_PG0_2_0_1680520037_0/m1_688_1652# INP COMP_PG0_2_0_1680520037_0/m1_1172_1316# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 COMP_PG0_2_0_1680520037_0/m1_1172_1316# INP COMP_PG0_2_0_1680520037_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 COMP_PG0_2_0_1680520037_0/m1_688_1652# VREF1 COMP_PG0_2_0_1680520037_0/li_749_1495# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X29 COMP_PG0_2_0_1680520037_0/li_749_1495# VREF1 COMP_PG0_2_0_1680520037_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X30 COMP_PG0_2_0_1680520037_0/m1_688_1652# VREF1 COMP_PG0_2_0_1680520037_0/li_749_1495# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 COMP_PG0_2_0_1680520037_0/li_749_1495# VREF1 COMP_PG0_2_0_1680520037_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X32 GND BIAS COMP_PG0_2_0_1680520037_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 COMP_PG0_2_0_1680520037_0/m1_688_1652# BIAS GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X34 GND BIAS COMP_PG0_2_0_1680520037_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X35 COMP_PG0_2_0_1680520037_0/m1_688_1652# BIAS GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X36 VCC COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/li_749_1495# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X37 COMP_PG0_2_0_1680520037_0/m1_1172_1316# COMP_PG0_2_0_1680520037_0/li_749_1495# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X38 COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/li_749_1495# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X39 VCC COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/li_749_1495# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X40 VCC COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/m1_1172_1316# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X41 COMP_PG0_2_0_1680520037_0/m1_1172_1316# COMP_PG0_2_0_1680520037_0/li_749_1495# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X42 COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/li_749_1495# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X43 VCC COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/m1_1172_1316# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X44 COMP_PG0_0_0_1680520035_0/m1_688_1652# VREF3 COMP_PG0_0_0_1680520035_0/m1_602_1568# GND sky130_fd_pr__nfet_01v8 ad=1.8312e+12p pd=1.78e+07u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X45 COMP_PG0_0_0_1680520035_0/m1_602_1568# VREF3 COMP_PG0_0_0_1680520035_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X46 COMP_PG0_0_0_1680520035_0/m1_688_1652# VREF3 COMP_PG0_0_0_1680520035_0/m1_602_1568# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X47 COMP_PG0_0_0_1680520035_0/m1_602_1568# VREF3 COMP_PG0_0_0_1680520035_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X48 COMP_PG0_0_0_1680520035_0/m1_688_1652# INP COMP_PG0_0_0_1680520035_0/m1_1172_1316# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X49 COMP_PG0_0_0_1680520035_0/m1_1172_1316# INP COMP_PG0_0_0_1680520035_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X50 COMP_PG0_0_0_1680520035_0/m1_688_1652# INP COMP_PG0_0_0_1680520035_0/m1_1172_1316# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X51 COMP_PG0_0_0_1680520035_0/m1_1172_1316# INP COMP_PG0_0_0_1680520035_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X52 GND COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X53 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_1172_1316# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X54 GND COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X55 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_1172_1316# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X56 GND COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_2720_1484# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X57 COMP_PG0_0_0_1680520035_0/m1_2720_1484# COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X58 GND COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_2720_1484# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X59 COMP_PG0_0_0_1680520035_0/m1_2720_1484# COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X60 COMP_PG0_0_0_1680520035_0/m1_2720_1484# COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X61 VCC COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_2720_1484# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X62 COMP_PG0_0_0_1680520035_0/m1_2720_1484# COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X63 VCC COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_2720_1484# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X64 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_1172_1316# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X65 VCC COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X66 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_1172_1316# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X67 VCC COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X68 GND BIAS COMP_PG0_0_0_1680520035_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X69 COMP_PG0_0_0_1680520035_0/m1_688_1652# BIAS GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X70 GND BIAS COMP_PG0_0_0_1680520035_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X71 COMP_PG0_0_0_1680520035_0/m1_688_1652# BIAS GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X72 VCC COMP_PG0_0_0_1680520035_0/m1_602_1568# COMP_PG0_0_0_1680520035_0/m1_602_1568# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X73 COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/m1_602_1568# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X74 COMP_PG0_0_0_1680520035_0/m1_602_1568# COMP_PG0_0_0_1680520035_0/m1_602_1568# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X75 VCC COMP_PG0_0_0_1680520035_0/m1_602_1568# COMP_PG0_0_0_1680520035_0/m1_602_1568# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X76 VCC COMP_PG0_0_0_1680520035_0/m1_602_1568# COMP_PG0_0_0_1680520035_0/m1_1172_1316# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X77 COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/m1_602_1568# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X78 COMP_PG0_0_0_1680520035_0/m1_602_1568# COMP_PG0_0_0_1680520035_0/m1_602_1568# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X79 VCC COMP_PG0_0_0_1680520035_0/m1_602_1568# COMP_PG0_0_0_1680520035_0/m1_1172_1316# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X80 C3 COMP_PG0_0_0_1680520035_0/m1_2720_1484# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X81 VCC COMP_PG0_0_0_1680520035_0/m1_2720_1484# C3 VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X82 C3 COMP_PG0_0_0_1680520035_0/m1_2720_1484# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X83 VCC COMP_PG0_0_0_1680520035_0/m1_2720_1484# C3 VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X84 GND COMP_PG0_0_0_1680520035_0/m1_2720_1484# C3 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X85 C3 COMP_PG0_0_0_1680520035_0/m1_2720_1484# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X86 GND COMP_PG0_0_0_1680520035_0/m1_2720_1484# C3 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X87 C3 COMP_PG0_0_0_1680520035_0/m1_2720_1484# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X88 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X89 VCC COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# COMP_PG0_1_0_1680520036_0/m1_2720_1484# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X90 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X91 VCC COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# COMP_PG0_1_0_1680520036_0/m1_2720_1484# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X92 COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# COMP_PG0_1_0_1680520036_0/m1_1172_1316# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X93 VCC COMP_PG0_1_0_1680520036_0/m1_1172_1316# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X94 COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# COMP_PG0_1_0_1680520036_0/m1_1172_1316# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X95 VCC COMP_PG0_1_0_1680520036_0/m1_1172_1316# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X96 GND COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# COMP_PG0_1_0_1680520036_0/m1_2720_1484# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X97 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X98 GND COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# COMP_PG0_1_0_1680520036_0/m1_2720_1484# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X99 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X100 GND COMP_PG0_1_0_1680520036_0/m1_1172_1316# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X101 COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# COMP_PG0_1_0_1680520036_0/m1_1172_1316# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X102 GND COMP_PG0_1_0_1680520036_0/m1_1172_1316# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X103 COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# COMP_PG0_1_0_1680520036_0/m1_1172_1316# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X104 COMP_PG0_1_0_1680520036_0/m1_688_1652# INP COMP_PG0_1_0_1680520036_0/m1_1172_1316# GND sky130_fd_pr__nfet_01v8 ad=1.8312e+12p pd=1.78e+07u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X105 COMP_PG0_1_0_1680520036_0/m1_1172_1316# INP COMP_PG0_1_0_1680520036_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X106 COMP_PG0_1_0_1680520036_0/m1_688_1652# INP COMP_PG0_1_0_1680520036_0/m1_1172_1316# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X107 COMP_PG0_1_0_1680520036_0/m1_1172_1316# INP COMP_PG0_1_0_1680520036_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X108 COMP_PG0_1_0_1680520036_0/m1_688_1652# VREF2 COMP_PG0_1_0_1680520036_0/m1_602_1568# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X109 COMP_PG0_1_0_1680520036_0/m1_602_1568# VREF2 COMP_PG0_1_0_1680520036_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X110 COMP_PG0_1_0_1680520036_0/m1_688_1652# VREF2 COMP_PG0_1_0_1680520036_0/m1_602_1568# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X111 COMP_PG0_1_0_1680520036_0/m1_602_1568# VREF2 COMP_PG0_1_0_1680520036_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X112 GND BIAS COMP_PG0_1_0_1680520036_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X113 COMP_PG0_1_0_1680520036_0/m1_688_1652# BIAS GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X114 GND BIAS COMP_PG0_1_0_1680520036_0/m1_688_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X115 COMP_PG0_1_0_1680520036_0/m1_688_1652# BIAS GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X116 VCC COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/m1_602_1568# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X117 COMP_PG0_1_0_1680520036_0/m1_1172_1316# COMP_PG0_1_0_1680520036_0/m1_602_1568# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X118 COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/m1_602_1568# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X119 VCC COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/m1_602_1568# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X120 VCC COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/m1_1172_1316# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X121 COMP_PG0_1_0_1680520036_0/m1_1172_1316# COMP_PG0_1_0_1680520036_0/m1_602_1568# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X122 COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/m1_602_1568# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X123 VCC COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/m1_1172_1316# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X124 C2 COMP_PG0_1_0_1680520036_0/m1_2720_1484# VCC VCC sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X125 VCC COMP_PG0_1_0_1680520036_0/m1_2720_1484# C2 VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X126 C2 COMP_PG0_1_0_1680520036_0/m1_2720_1484# VCC VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X127 VCC COMP_PG0_1_0_1680520036_0/m1_2720_1484# C2 VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X128 GND COMP_PG0_1_0_1680520036_0/m1_2720_1484# C2 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X129 C2 COMP_PG0_1_0_1680520036_0/m1_2720_1484# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X130 GND COMP_PG0_1_0_1680520036_0/m1_2720_1484# C2 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X131 C2 COMP_PG0_1_0_1680520036_0/m1_2720_1484# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.59fF
C1 COMP_PG0_0_0_1680520035_0/m1_602_1568# COMP_PG0_0_0_1680520035_0/m1_2720_1484# 0.00fF
C2 VREF3 BIAS 0.00fF
C3 COMP_PG0_1_0_1680520036_0/m1_602_1568# INP 0.01fF
C4 COMP_PG0_0_0_1680520035_0/m1_602_1568# C2 0.00fF
C5 VREF3 INP 0.31fF
C6 COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/m1_688_1652# 1.72fF
C7 VREF1 VCC 0.03fF
C8 BIAS COMP_PG0_2_0_1680520037_0/m1_1172_1316# 0.00fF
C9 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_688_1652# 0.00fF
C10 C3 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# 0.00fF
C11 COMP_PG0_2_0_1680520037_0/m1_2720_1484# INP 0.00fF
C12 INP COMP_PG0_2_0_1680520037_0/m1_1172_1316# 0.26fF
C13 VREF1 COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.24fF
C14 VREF3 COMP_PG0_0_0_1680520035_0/m1_602_1568# 0.22fF
C15 COMP_PG0_1_0_1680520036_0/m1_688_1652# COMP_PG0_2_0_1680520037_0/m1_1172_1316# 0.00fF
C16 COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# 0.01fF
C17 COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_2_0_1680520037_0/li_749_1495# 0.00fF
C18 VCC VREF2 0.06fF
C19 VREF2 COMP_PG0_1_0_1680520036_0/m1_1172_1316# 0.00fF
C20 VCC BIAS 1.24fF
C21 VREF2 COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.00fF
C22 INP VCC 5.30fF
C23 BIAS COMP_PG0_1_0_1680520036_0/m1_1172_1316# 0.47fF
C24 COMP_PG0_2_0_1680520037_0/m1_2720_1484# COMP_PG0_2_0_1680520037_0/li_749_1495# 0.00fF
C25 COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/m1_1172_1316# 0.94fF
C26 BIAS COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.22fF
C27 INP COMP_PG0_1_0_1680520036_0/m1_1172_1316# 0.56fF
C28 COMP_PG0_1_0_1680520036_0/m1_688_1652# VCC 0.40fF
C29 COMP_PG0_0_0_1680520035_0/m1_1172_1316# BIAS 0.00fF
C30 INP COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.27fF
C31 COMP_PG0_2_0_1680520037_0/m1_2720_1484# COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# 0.60fF
C32 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_1172_1316# 1.01fF
C33 COMP_PG0_1_0_1680520036_0/m1_688_1652# COMP_PG0_1_0_1680520036_0/m1_1172_1316# 1.38fF
C34 COMP_PG0_0_0_1680520035_0/m1_1172_1316# INP 0.26fF
C35 VCC COMP_PG0_0_0_1680520035_0/m1_602_1568# 4.64fF
C36 COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_2_0_1680520037_0/m1_1172_1316# 0.00fF
C37 COMP_PG0_1_0_1680520036_0/m1_688_1652# COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.06fF
C38 VCC COMP_PG0_0_0_1680520035_0/m1_2720_1484# 3.75fF
C39 COMP_PG0_2_0_1680520037_0/li_749_1495# VCC 4.67fF
C40 COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/m1_602_1568# 1.08fF
C41 VCC C2 1.63fF
C42 COMP_PG0_2_0_1680520037_0/m1_2720_1484# COMP_PG0_2_0_1680520037_0/m1_1172_1316# 0.01fF
C43 VREF2 COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.00fF
C44 COMP_PG0_0_0_1680520035_0/m1_688_1652# BIAS 0.22fF
C45 COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_1_0_1680520036_0/m1_1172_1316# 0.00fF
C46 COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/m1_2720_1484# 0.01fF
C47 C2 COMP_PG0_1_0_1680520036_0/m1_1172_1316# 0.00fF
C48 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# VCC 4.34fF
C49 INP COMP_PG0_0_0_1680520035_0/m1_688_1652# 0.28fF
C50 COMP_PG0_2_0_1680520037_0/li_749_1495# COMP_PG0_2_0_1680520037_0/m1_688_1652# 1.65fF
C51 BIAS COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.71fF
C52 COMP_PG0_1_0_1680520036_0/m1_602_1568# VCC 4.72fF
C53 COMP_PG0_0_0_1680520035_0/m1_1172_1316# C2 0.00fF
C54 INP COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.49fF
C55 VREF3 VCC 0.04fF
C56 COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/m1_1172_1316# 1.05fF
C57 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.00fF
C58 COMP_PG0_1_0_1680520036_0/m1_688_1652# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.00fF
C59 COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.00fF
C60 COMP_PG0_0_0_1680520035_0/m1_688_1652# COMP_PG0_0_0_1680520035_0/m1_602_1568# 1.72fF
C61 COMP_PG0_2_0_1680520037_0/m1_2720_1484# VCC 3.79fF
C62 COMP_PG0_1_0_1680520036_0/m1_2720_1484# BIAS 0.59fF
C63 VCC COMP_PG0_2_0_1680520037_0/m1_1172_1316# 4.43fF
C64 VREF3 COMP_PG0_0_0_1680520035_0/m1_1172_1316# 0.00fF
C65 COMP_PG0_0_0_1680520035_0/m1_688_1652# COMP_PG0_0_0_1680520035_0/m1_2720_1484# 0.00fF
C66 C3 COMP_PG0_0_0_1680520035_0/m1_2720_1484# 0.78fF
C67 COMP_PG0_1_0_1680520036_0/m1_2720_1484# INP 0.30fF
C68 COMP_PG0_0_0_1680520035_0/m1_688_1652# C2 0.02fF
C69 COMP_PG0_2_0_1680520037_0/m1_2720_1484# COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.00fF
C70 COMP_PG0_2_0_1680520037_0/m1_1172_1316# COMP_PG0_2_0_1680520037_0/m1_688_1652# 1.34fF
C71 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_1_0_1680520036_0/m1_688_1652# 0.00fF
C72 C2 COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.00fF
C73 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_0_0_1680520035_0/m1_602_1568# 0.00fF
C74 VREF3 COMP_PG0_0_0_1680520035_0/m1_688_1652# 0.24fF
C75 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# INP 0.00fF
C76 COMP_PG0_1_0_1680520036_0/m1_602_1568# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.01fF
C77 C1 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# 0.00fF
C78 VCC COMP_PG0_1_0_1680520036_0/m1_1172_1316# 4.16fF
C79 VREF3 COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.00fF
C80 COMP_PG0_1_0_1680520036_0/m1_2720_1484# C2 0.76fF
C81 VCC COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.26fF
C82 COMP_PG0_0_0_1680520035_0/m1_1172_1316# VCC 4.37fF
C83 COMP_PG0_1_0_1680520036_0/m1_1172_1316# COMP_PG0_2_0_1680520037_0/m1_688_1652# 0.00fF
C84 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_602_1568# 0.01fF
C85 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_1_0_1680520036_0/m1_602_1568# 0.00fF
C86 VREF1 VREF2 0.02fF
C87 C1 COMP_PG0_2_0_1680520037_0/m1_2720_1484# 0.77fF
C88 C1 COMP_PG0_2_0_1680520037_0/m1_1172_1316# 0.00fF
C89 COMP_PG0_1_0_1680520036_0/m1_2720_1484# VREF3 0.03fF
C90 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_2720_1484# 0.60fF
C91 VREF1 BIAS 0.00fF
C92 INP VREF1 0.33fF
C93 VCC COMP_PG0_0_0_1680520035_0/m1_688_1652# 0.37fF
C94 C3 VCC 1.63fF
C95 COMP_PG0_1_0_1680520036_0/m1_688_1652# VREF1 0.00fF
C96 VCC COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 4.15fF
C97 VREF3 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# 0.00fF
C98 C1 VCC 1.65fF
C99 C3 COMP_PG0_0_0_1680520035_0/m1_1172_1316# 0.00fF
C100 COMP_PG0_0_0_1680520035_0/m1_1172_1316# COMP_PG0_0_0_1680520035_0/m1_688_1652# 1.38fF
C101 VREF2 BIAS 0.00fF
C102 COMP_PG0_1_0_1680520036_0/m1_1172_1316# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 1.01fF
C103 INP VREF2 0.31fF
C104 COMP_PG0_1_0_1680520036_0/m1_2720_1484# VCC 3.67fF
C105 COMP_PG0_1_0_1680520036_0/m1_688_1652# VREF2 0.24fF
C106 COMP_PG0_2_0_1680520037_0/li_749_1495# VREF1 0.22fF
C107 INP BIAS 0.00fF
C108 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_1_0_1680520036_0/m1_1172_1316# 0.01fF
C109 COMP_PG0_1_0_1680520036_0/m1_688_1652# BIAS 0.23fF
C110 VREF1 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# 0.00fF
C111 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_0_0_1680520035_0/m1_1172_1316# 0.00fF
C112 COMP_PG0_1_0_1680520036_0/m1_688_1652# INP 0.28fF
C113 COMP_PG0_0_0_1680520035_0/m1_602_1568# BIAS 0.04fF
C114 COMP_PG0_0_0_1680520035_0/m1_688_1652# COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# 0.00fF
C115 INP COMP_PG0_0_0_1680520035_0/m1_602_1568# 0.01fF
C116 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# VCC 4.43fF
C117 COMP_PG0_2_0_1680520037_0/li_749_1495# BIAS 0.04fF
C118 INP COMP_PG0_0_0_1680520035_0/m1_2720_1484# 0.00fF
C119 C2 BIAS 0.04fF
C120 VREF1 COMP_PG0_2_0_1680520037_0/m1_1172_1316# 0.00fF
C121 COMP_PG0_2_0_1680520037_0/li_749_1495# INP 0.01fF
C122 COMP_PG0_1_0_1680520036_0/m1_602_1568# VREF2 0.22fF
C123 INP C2 0.00fF
C124 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# COMP_PG0_0_0_1680520035_0/m1_1172_1316# 1.02fF
C125 COMP_PG0_1_0_1680520036_0/m1_2720_1484# COMP_PG0_0_0_1680520035_0/m1_688_1652# 0.01fF
C126 COMP_PG0_1_0_1680520036_0/m1_688_1652# COMP_PG0_2_0_1680520037_0/li_749_1495# 0.00fF
C127 COMP_PG0_1_0_1680520036_0/m1_602_1568# BIAS 0.92fF
C128 INP COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# 0.00fF
C129 BIAS GND 1.97fF
C130 C2 GND 1.32fF
C131 COMP_PG0_1_0_1680520036_0/m1_602_1568# GND 0.37fF
C132 VREF2 GND 1.25fF
C133 COMP_PG0_1_0_1680520036_0/m1_688_1652# GND 1.89fF
C134 COMP_PG0_1_0_1680520036_0/m1_1172_1316# GND 1.35fF
C135 COMP_PG0_1_0_1680520036_0/m1_2720_1484# GND 2.81fF
C136 COMP_PG0_1_0_1680520036_0/STAGE2_INV_90501218_PG0_1_0_1680520031_1680520036_0/li_663_571# GND 1.97fF
C137 C3 GND 1.38fF
C138 COMP_PG0_0_0_1680520035_0/m1_1172_1316# GND 1.46fF
C139 COMP_PG0_0_0_1680520035_0/m1_2720_1484# GND 2.71fF
C140 COMP_PG0_0_0_1680520035_0/STAGE2_INV_90501218_PG0_0_0_1680520030_1680520035_0/li_663_571# GND 2.05fF
C141 COMP_PG0_0_0_1680520035_0/m1_688_1652# GND 1.84fF
C142 COMP_PG0_0_0_1680520035_0/m1_602_1568# GND 0.35fF
C143 VREF3 GND 1.24fF
C144 COMP_PG0_2_0_1680520037_0/m1_1172_1316# GND 1.54fF
C145 COMP_PG0_2_0_1680520037_0/li_749_1495# GND 0.10fF
C146 VREF1 GND 1.18fF
C147 COMP_PG0_2_0_1680520037_0/m1_688_1652# GND 1.97fF
C148 VCC GND 50.25fF
C149 COMP_PG0_2_0_1680520037_0/m1_2720_1484# GND 2.76fF
C150 COMP_PG0_2_0_1680520037_0/STAGE2_INV_90501218_PG0_2_0_1680520031_1680520037_0/li_663_571# GND 2.09fF
C151 C1 GND 1.35fF
.ends TWOBIT_FLASH_ADC

x1 GND VCC C3 C2 C1 VREF2 VREF3 VREF1 BIAS INP TWOBIT_FLASH_ADC
V1 VCC GND 3.3
V2 BIAS GND 0.9
V3 VREF1 GND 0.7
V4 VREF2 GND 1.4
V5 VREF3 GND 2.1
V6 INP GND sine(0 3.3 600000000)

.tran 10p 20n
.control
run
plot v(VREF1) v(VREF2) v(VREF3) v(INP) v(C3) v(C2) v(C1)
save all
.endc

