MACRO TWOBIT_FLASH_ADC
  ORIGIN 0 0 ;
  FOREIGN TWOBIT_FLASH_ADC 0 0 ;
  SIZE 57.35 BY 15.71 ;
  PIN BIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.6 12.04 17.8 12.32 ;
      LAYER M2 ;
        RECT 20.04 12.04 21.24 12.32 ;
      LAYER M2 ;
        RECT 38.96 12.04 40.16 12.32 ;
      LAYER M2 ;
        RECT 17.63 12.04 20.21 12.32 ;
      LAYER M2 ;
        RECT 21.07 12.04 22.79 12.32 ;
      LAYER M1 ;
        RECT 22.665 11.76 22.915 12.18 ;
      LAYER M2 ;
        RECT 22.79 11.62 37.41 11.9 ;
      LAYER M1 ;
        RECT 37.285 11.76 37.535 12.18 ;
      LAYER M2 ;
        RECT 37.41 12.04 39.13 12.32 ;
    END
  END BIAS
  PIN VREF3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 39.82 2.8 41.02 3.08 ;
    END
  END VREF3
  PIN INP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
      LAYER M2 ;
        RECT 24.34 2.8 25.54 3.08 ;
      LAYER M2 ;
        RECT 43.26 2.8 44.46 3.08 ;
      LAYER M2 ;
        RECT 13.33 2.8 15.05 3.08 ;
      LAYER M1 ;
        RECT 14.925 2.52 15.175 2.94 ;
      LAYER M2 ;
        RECT 15.05 2.38 24.51 2.66 ;
      LAYER M3 ;
        RECT 24.37 2.52 24.65 2.94 ;
      LAYER M2 ;
        RECT 24.35 2.8 24.67 3.08 ;
      LAYER M2 ;
        RECT 24.51 2.38 43 2.66 ;
      LAYER M1 ;
        RECT 42.875 2.52 43.125 2.94 ;
      LAYER M2 ;
        RECT 43 2.8 43.43 3.08 ;
    END
  END INP
  PIN C3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 54.44 7 55.64 7.28 ;
      LAYER M2 ;
        RECT 54.44 7.84 55.64 8.12 ;
      LAYER M2 ;
        RECT 54.88 7 55.2 7.28 ;
      LAYER M3 ;
        RECT 54.9 7.14 55.18 7.98 ;
      LAYER M2 ;
        RECT 54.88 7.84 55.2 8.12 ;
    END
  END C3
  PIN VREF2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 20.9 2.8 22.1 3.08 ;
    END
  END VREF2
  PIN C2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 35.52 7 36.72 7.28 ;
      LAYER M2 ;
        RECT 35.52 7.84 36.72 8.12 ;
      LAYER M2 ;
        RECT 35.96 7 36.28 7.28 ;
      LAYER M3 ;
        RECT 35.98 7.14 36.26 7.98 ;
      LAYER M2 ;
        RECT 35.96 7.84 36.28 8.12 ;
    END
  END C2
  PIN VREF1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 15.74 2.8 16.94 3.08 ;
    END
  END VREF1
  PIN C1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
      LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
      LAYER M2 ;
        RECT 1.56 7 1.88 7.28 ;
      LAYER M3 ;
        RECT 1.58 7.14 1.86 7.98 ;
      LAYER M2 ;
        RECT 1.56 7.84 1.88 8.12 ;
    END
  END C1
  OBS 
  LAYER M2 ;
        RECT 43.26 7 44.46 7.28 ;
  LAYER M2 ;
        RECT 43.26 8.26 44.46 8.54 ;
  LAYER M2 ;
        RECT 47.56 2.8 48.76 3.08 ;
  LAYER M2 ;
        RECT 47.56 12.04 48.76 12.32 ;
  LAYER M2 ;
        RECT 48 2.8 48.32 3.08 ;
  LAYER M3 ;
        RECT 48.02 2.94 48.3 12.18 ;
  LAYER M2 ;
        RECT 48 12.04 48.32 12.32 ;
  LAYER M2 ;
        RECT 43.7 7 44.02 7.28 ;
  LAYER M3 ;
        RECT 43.72 7.14 44 8.4 ;
  LAYER M2 ;
        RECT 43.7 8.26 44.02 8.54 ;
  LAYER M3 ;
        RECT 43.72 7.375 44 7.745 ;
  LAYER M2 ;
        RECT 43.86 7.42 48.16 7.7 ;
  LAYER M3 ;
        RECT 48.02 7.375 48.3 7.745 ;
  LAYER M2 ;
        RECT 43.7 7 44.02 7.28 ;
  LAYER M3 ;
        RECT 43.72 6.98 44 7.3 ;
  LAYER M2 ;
        RECT 43.7 8.26 44.02 8.54 ;
  LAYER M3 ;
        RECT 43.72 8.24 44 8.56 ;
  LAYER M2 ;
        RECT 43.7 7 44.02 7.28 ;
  LAYER M3 ;
        RECT 43.72 6.98 44 7.3 ;
  LAYER M2 ;
        RECT 43.7 8.26 44.02 8.54 ;
  LAYER M3 ;
        RECT 43.72 8.24 44 8.56 ;
  LAYER M2 ;
        RECT 43.7 7 44.02 7.28 ;
  LAYER M3 ;
        RECT 43.72 6.98 44 7.3 ;
  LAYER M2 ;
        RECT 43.7 7.42 44.02 7.7 ;
  LAYER M3 ;
        RECT 43.72 7.4 44 7.72 ;
  LAYER M2 ;
        RECT 43.7 8.26 44.02 8.54 ;
  LAYER M3 ;
        RECT 43.72 8.24 44 8.56 ;
  LAYER M2 ;
        RECT 48 7.42 48.32 7.7 ;
  LAYER M3 ;
        RECT 48.02 7.4 48.3 7.72 ;
  LAYER M2 ;
        RECT 43.7 7 44.02 7.28 ;
  LAYER M3 ;
        RECT 43.72 6.98 44 7.3 ;
  LAYER M2 ;
        RECT 43.7 7.42 44.02 7.7 ;
  LAYER M3 ;
        RECT 43.72 7.4 44 7.72 ;
  LAYER M2 ;
        RECT 43.7 8.26 44.02 8.54 ;
  LAYER M3 ;
        RECT 43.72 8.24 44 8.56 ;
  LAYER M2 ;
        RECT 48 7.42 48.32 7.7 ;
  LAYER M3 ;
        RECT 48.02 7.4 48.3 7.72 ;
  LAYER M2 ;
        RECT 54.44 2.8 55.64 3.08 ;
  LAYER M2 ;
        RECT 54.44 12.04 55.64 12.32 ;
  LAYER M2 ;
        RECT 54.45 2.8 54.77 3.08 ;
  LAYER M3 ;
        RECT 54.47 2.94 54.75 12.18 ;
  LAYER M2 ;
        RECT 54.45 12.04 54.77 12.32 ;
  LAYER M2 ;
        RECT 51 7 52.2 7.28 ;
  LAYER M2 ;
        RECT 51 7.84 52.2 8.12 ;
  LAYER M2 ;
        RECT 51.44 7 51.76 7.28 ;
  LAYER M3 ;
        RECT 51.46 7.14 51.74 7.98 ;
  LAYER M2 ;
        RECT 51.44 7.84 51.76 8.12 ;
  LAYER M3 ;
        RECT 54.47 7.375 54.75 7.745 ;
  LAYER M2 ;
        RECT 51.6 7.42 54.61 7.7 ;
  LAYER M3 ;
        RECT 51.46 7.375 51.74 7.745 ;
  LAYER M2 ;
        RECT 51.44 7.42 51.76 7.7 ;
  LAYER M3 ;
        RECT 51.46 7.4 51.74 7.72 ;
  LAYER M2 ;
        RECT 54.45 7.42 54.77 7.7 ;
  LAYER M3 ;
        RECT 54.47 7.4 54.75 7.72 ;
  LAYER M2 ;
        RECT 51.44 7.42 51.76 7.7 ;
  LAYER M3 ;
        RECT 51.46 7.4 51.74 7.72 ;
  LAYER M2 ;
        RECT 54.45 7.42 54.77 7.7 ;
  LAYER M3 ;
        RECT 54.47 7.4 54.75 7.72 ;
  LAYER M2 ;
        RECT 39.82 7 41.02 7.28 ;
  LAYER M3 ;
        RECT 43.29 7.82 43.57 12.34 ;
  LAYER M2 ;
        RECT 40.85 7 42.57 7.28 ;
  LAYER M3 ;
        RECT 42.43 7.14 42.71 7.56 ;
  LAYER M4 ;
        RECT 42.57 7.16 43.43 7.96 ;
  LAYER M3 ;
        RECT 43.29 7.56 43.57 7.98 ;
  LAYER M2 ;
        RECT 42.41 7 42.73 7.28 ;
  LAYER M3 ;
        RECT 42.43 6.98 42.71 7.3 ;
  LAYER M3 ;
        RECT 42.43 7.375 42.71 7.745 ;
  LAYER M4 ;
        RECT 42.405 7.16 42.735 7.96 ;
  LAYER M3 ;
        RECT 43.29 7.375 43.57 7.745 ;
  LAYER M4 ;
        RECT 43.265 7.16 43.595 7.96 ;
  LAYER M2 ;
        RECT 42.41 7 42.73 7.28 ;
  LAYER M3 ;
        RECT 42.43 6.98 42.71 7.3 ;
  LAYER M3 ;
        RECT 42.43 7.375 42.71 7.745 ;
  LAYER M4 ;
        RECT 42.405 7.16 42.735 7.96 ;
  LAYER M3 ;
        RECT 43.29 7.375 43.57 7.745 ;
  LAYER M4 ;
        RECT 43.265 7.16 43.595 7.96 ;
  LAYER M2 ;
        RECT 39.39 6.58 41.45 6.86 ;
  LAYER M2 ;
        RECT 38.96 7.84 40.16 8.12 ;
  LAYER M2 ;
        RECT 42.83 6.58 44.89 6.86 ;
  LAYER M2 ;
        RECT 39.4 6.58 39.72 6.86 ;
  LAYER M3 ;
        RECT 39.42 6.72 39.7 7.98 ;
  LAYER M2 ;
        RECT 39.4 7.84 39.72 8.12 ;
  LAYER M2 ;
        RECT 41.28 6.58 43 6.86 ;
  LAYER M2 ;
        RECT 39.4 6.58 39.72 6.86 ;
  LAYER M3 ;
        RECT 39.42 6.56 39.7 6.88 ;
  LAYER M2 ;
        RECT 39.4 7.84 39.72 8.12 ;
  LAYER M3 ;
        RECT 39.42 7.82 39.7 8.14 ;
  LAYER M2 ;
        RECT 39.4 6.58 39.72 6.86 ;
  LAYER M3 ;
        RECT 39.42 6.56 39.7 6.88 ;
  LAYER M2 ;
        RECT 39.4 7.84 39.72 8.12 ;
  LAYER M3 ;
        RECT 39.42 7.82 39.7 8.14 ;
  LAYER M2 ;
        RECT 39.4 6.58 39.72 6.86 ;
  LAYER M3 ;
        RECT 39.42 6.56 39.7 6.88 ;
  LAYER M2 ;
        RECT 39.4 7.84 39.72 8.12 ;
  LAYER M3 ;
        RECT 39.42 7.82 39.7 8.14 ;
  LAYER M2 ;
        RECT 39.4 6.58 39.72 6.86 ;
  LAYER M3 ;
        RECT 39.42 6.56 39.7 6.88 ;
  LAYER M2 ;
        RECT 39.4 7.84 39.72 8.12 ;
  LAYER M3 ;
        RECT 39.42 7.82 39.7 8.14 ;
  LAYER M2 ;
        RECT 51 2.8 52.2 3.08 ;
  LAYER M2 ;
        RECT 47.56 7 48.76 7.28 ;
  LAYER M2 ;
        RECT 47.56 7.84 48.76 8.12 ;
  LAYER M2 ;
        RECT 51 12.04 52.2 12.32 ;
  LAYER M2 ;
        RECT 49.88 2.8 51.17 3.08 ;
  LAYER M1 ;
        RECT 49.755 2.94 50.005 7.14 ;
  LAYER M2 ;
        RECT 48.59 7 49.88 7.28 ;
  LAYER M2 ;
        RECT 48.43 7 48.75 7.28 ;
  LAYER M3 ;
        RECT 48.45 7.14 48.73 7.98 ;
  LAYER M2 ;
        RECT 48.43 7.84 48.75 8.12 ;
  LAYER M1 ;
        RECT 49.755 7.14 50.005 12.18 ;
  LAYER M2 ;
        RECT 49.88 12.04 51.17 12.32 ;
  LAYER M1 ;
        RECT 49.755 2.855 50.005 3.025 ;
  LAYER M2 ;
        RECT 49.71 2.8 50.05 3.08 ;
  LAYER M1 ;
        RECT 49.755 7.055 50.005 7.225 ;
  LAYER M2 ;
        RECT 49.71 7 50.05 7.28 ;
  LAYER M1 ;
        RECT 49.755 2.855 50.005 3.025 ;
  LAYER M2 ;
        RECT 49.71 2.8 50.05 3.08 ;
  LAYER M1 ;
        RECT 49.755 7.055 50.005 7.225 ;
  LAYER M2 ;
        RECT 49.71 7 50.05 7.28 ;
  LAYER M1 ;
        RECT 49.755 2.855 50.005 3.025 ;
  LAYER M2 ;
        RECT 49.71 2.8 50.05 3.08 ;
  LAYER M1 ;
        RECT 49.755 7.055 50.005 7.225 ;
  LAYER M2 ;
        RECT 49.71 7 50.05 7.28 ;
  LAYER M2 ;
        RECT 48.43 7 48.75 7.28 ;
  LAYER M3 ;
        RECT 48.45 6.98 48.73 7.3 ;
  LAYER M2 ;
        RECT 48.43 7.84 48.75 8.12 ;
  LAYER M3 ;
        RECT 48.45 7.82 48.73 8.14 ;
  LAYER M1 ;
        RECT 49.755 2.855 50.005 3.025 ;
  LAYER M2 ;
        RECT 49.71 2.8 50.05 3.08 ;
  LAYER M1 ;
        RECT 49.755 7.055 50.005 7.225 ;
  LAYER M2 ;
        RECT 49.71 7 50.05 7.28 ;
  LAYER M2 ;
        RECT 48.43 7 48.75 7.28 ;
  LAYER M3 ;
        RECT 48.45 6.98 48.73 7.3 ;
  LAYER M2 ;
        RECT 48.43 7.84 48.75 8.12 ;
  LAYER M3 ;
        RECT 48.45 7.82 48.73 8.14 ;
  LAYER M1 ;
        RECT 49.755 2.855 50.005 3.025 ;
  LAYER M2 ;
        RECT 49.71 2.8 50.05 3.08 ;
  LAYER M1 ;
        RECT 49.755 7.055 50.005 7.225 ;
  LAYER M2 ;
        RECT 49.71 7 50.05 7.28 ;
  LAYER M1 ;
        RECT 49.755 12.095 50.005 12.265 ;
  LAYER M2 ;
        RECT 49.71 12.04 50.05 12.32 ;
  LAYER M2 ;
        RECT 48.43 7 48.75 7.28 ;
  LAYER M3 ;
        RECT 48.45 6.98 48.73 7.3 ;
  LAYER M2 ;
        RECT 48.43 7.84 48.75 8.12 ;
  LAYER M3 ;
        RECT 48.45 7.82 48.73 8.14 ;
  LAYER M1 ;
        RECT 49.755 2.855 50.005 3.025 ;
  LAYER M2 ;
        RECT 49.71 2.8 50.05 3.08 ;
  LAYER M1 ;
        RECT 49.755 7.055 50.005 7.225 ;
  LAYER M2 ;
        RECT 49.71 7 50.05 7.28 ;
  LAYER M1 ;
        RECT 49.755 12.095 50.005 12.265 ;
  LAYER M2 ;
        RECT 49.71 12.04 50.05 12.32 ;
  LAYER M2 ;
        RECT 48.43 7 48.75 7.28 ;
  LAYER M3 ;
        RECT 48.45 6.98 48.73 7.3 ;
  LAYER M2 ;
        RECT 48.43 7.84 48.75 8.12 ;
  LAYER M3 ;
        RECT 48.45 7.82 48.73 8.14 ;
  LAYER M1 ;
        RECT 48.465 7.895 48.715 11.425 ;
  LAYER M1 ;
        RECT 48.465 11.675 48.715 12.685 ;
  LAYER M1 ;
        RECT 48.465 13.775 48.715 14.785 ;
  LAYER M1 ;
        RECT 48.895 7.895 49.145 11.425 ;
  LAYER M1 ;
        RECT 48.035 7.895 48.285 11.425 ;
  LAYER M1 ;
        RECT 47.605 7.895 47.855 11.425 ;
  LAYER M1 ;
        RECT 47.605 11.675 47.855 12.685 ;
  LAYER M1 ;
        RECT 47.605 13.775 47.855 14.785 ;
  LAYER M1 ;
        RECT 47.175 7.895 47.425 11.425 ;
  LAYER M2 ;
        RECT 47.56 14.14 48.76 14.42 ;
  LAYER M2 ;
        RECT 47.13 8.26 49.19 8.54 ;
  LAYER M2 ;
        RECT 47.56 7.84 48.76 8.12 ;
  LAYER M2 ;
        RECT 47.56 12.04 48.76 12.32 ;
  LAYER M3 ;
        RECT 47.59 8.24 47.87 14.44 ;
  LAYER M1 ;
        RECT 51.905 7.895 52.155 11.425 ;
  LAYER M1 ;
        RECT 51.905 11.675 52.155 12.685 ;
  LAYER M1 ;
        RECT 51.905 13.775 52.155 14.785 ;
  LAYER M1 ;
        RECT 52.335 7.895 52.585 11.425 ;
  LAYER M1 ;
        RECT 51.475 7.895 51.725 11.425 ;
  LAYER M1 ;
        RECT 51.045 7.895 51.295 11.425 ;
  LAYER M1 ;
        RECT 51.045 11.675 51.295 12.685 ;
  LAYER M1 ;
        RECT 51.045 13.775 51.295 14.785 ;
  LAYER M1 ;
        RECT 50.615 7.895 50.865 11.425 ;
  LAYER M2 ;
        RECT 51 14.14 52.2 14.42 ;
  LAYER M2 ;
        RECT 50.57 8.26 52.63 8.54 ;
  LAYER M2 ;
        RECT 51 7.84 52.2 8.12 ;
  LAYER M2 ;
        RECT 51 12.04 52.2 12.32 ;
  LAYER M3 ;
        RECT 51.03 8.24 51.31 14.44 ;
  LAYER M1 ;
        RECT 48.465 3.695 48.715 7.225 ;
  LAYER M1 ;
        RECT 48.465 2.435 48.715 3.445 ;
  LAYER M1 ;
        RECT 48.465 0.335 48.715 1.345 ;
  LAYER M1 ;
        RECT 48.895 3.695 49.145 7.225 ;
  LAYER M1 ;
        RECT 48.035 3.695 48.285 7.225 ;
  LAYER M1 ;
        RECT 47.605 3.695 47.855 7.225 ;
  LAYER M1 ;
        RECT 47.605 2.435 47.855 3.445 ;
  LAYER M1 ;
        RECT 47.605 0.335 47.855 1.345 ;
  LAYER M1 ;
        RECT 47.175 3.695 47.425 7.225 ;
  LAYER M2 ;
        RECT 47.56 0.7 48.76 0.98 ;
  LAYER M2 ;
        RECT 47.13 6.58 49.19 6.86 ;
  LAYER M2 ;
        RECT 47.56 7 48.76 7.28 ;
  LAYER M2 ;
        RECT 47.56 2.8 48.76 3.08 ;
  LAYER M3 ;
        RECT 47.59 0.68 47.87 6.88 ;
  LAYER M1 ;
        RECT 51.905 3.695 52.155 7.225 ;
  LAYER M1 ;
        RECT 51.905 2.435 52.155 3.445 ;
  LAYER M1 ;
        RECT 51.905 0.335 52.155 1.345 ;
  LAYER M1 ;
        RECT 52.335 3.695 52.585 7.225 ;
  LAYER M1 ;
        RECT 51.475 3.695 51.725 7.225 ;
  LAYER M1 ;
        RECT 51.045 3.695 51.295 7.225 ;
  LAYER M1 ;
        RECT 51.045 2.435 51.295 3.445 ;
  LAYER M1 ;
        RECT 51.045 0.335 51.295 1.345 ;
  LAYER M1 ;
        RECT 50.615 3.695 50.865 7.225 ;
  LAYER M2 ;
        RECT 51 0.7 52.2 0.98 ;
  LAYER M2 ;
        RECT 50.57 6.58 52.63 6.86 ;
  LAYER M2 ;
        RECT 51 7 52.2 7.28 ;
  LAYER M2 ;
        RECT 51 2.8 52.2 3.08 ;
  LAYER M3 ;
        RECT 51.03 0.68 51.31 6.88 ;
  LAYER M1 ;
        RECT 42.445 7.895 42.695 11.425 ;
  LAYER M1 ;
        RECT 42.445 11.675 42.695 12.685 ;
  LAYER M1 ;
        RECT 42.445 13.775 42.695 14.785 ;
  LAYER M1 ;
        RECT 42.015 7.895 42.265 11.425 ;
  LAYER M1 ;
        RECT 42.875 7.895 43.125 11.425 ;
  LAYER M1 ;
        RECT 43.305 7.895 43.555 11.425 ;
  LAYER M1 ;
        RECT 43.305 11.675 43.555 12.685 ;
  LAYER M1 ;
        RECT 43.305 13.775 43.555 14.785 ;
  LAYER M1 ;
        RECT 43.735 7.895 43.985 11.425 ;
  LAYER M1 ;
        RECT 44.165 7.895 44.415 11.425 ;
  LAYER M1 ;
        RECT 44.165 11.675 44.415 12.685 ;
  LAYER M1 ;
        RECT 44.165 13.775 44.415 14.785 ;
  LAYER M1 ;
        RECT 44.595 7.895 44.845 11.425 ;
  LAYER M1 ;
        RECT 45.025 7.895 45.275 11.425 ;
  LAYER M1 ;
        RECT 45.025 11.675 45.275 12.685 ;
  LAYER M1 ;
        RECT 45.025 13.775 45.275 14.785 ;
  LAYER M1 ;
        RECT 45.455 7.895 45.705 11.425 ;
  LAYER M2 ;
        RECT 42.4 12.04 45.32 12.32 ;
  LAYER M2 ;
        RECT 42.4 7.84 45.32 8.12 ;
  LAYER M2 ;
        RECT 42.4 14.14 45.32 14.42 ;
  LAYER M2 ;
        RECT 41.97 8.68 45.75 8.96 ;
  LAYER M3 ;
        RECT 43.29 7.82 43.57 12.34 ;
  LAYER M2 ;
        RECT 43.26 8.26 44.46 8.54 ;
  LAYER M3 ;
        RECT 44.15 8.66 44.43 14.44 ;
  LAYER M1 ;
        RECT 54.485 7.895 54.735 11.425 ;
  LAYER M1 ;
        RECT 54.485 11.675 54.735 12.685 ;
  LAYER M1 ;
        RECT 54.485 13.775 54.735 14.785 ;
  LAYER M1 ;
        RECT 54.055 7.895 54.305 11.425 ;
  LAYER M1 ;
        RECT 54.915 7.895 55.165 11.425 ;
  LAYER M1 ;
        RECT 55.345 7.895 55.595 11.425 ;
  LAYER M1 ;
        RECT 55.345 11.675 55.595 12.685 ;
  LAYER M1 ;
        RECT 55.345 13.775 55.595 14.785 ;
  LAYER M1 ;
        RECT 55.775 7.895 56.025 11.425 ;
  LAYER M2 ;
        RECT 54.44 14.14 55.64 14.42 ;
  LAYER M2 ;
        RECT 54.01 8.26 56.07 8.54 ;
  LAYER M2 ;
        RECT 54.44 7.84 55.64 8.12 ;
  LAYER M2 ;
        RECT 54.44 12.04 55.64 12.32 ;
  LAYER M3 ;
        RECT 55.33 8.24 55.61 14.44 ;
  LAYER M1 ;
        RECT 54.485 3.695 54.735 7.225 ;
  LAYER M1 ;
        RECT 54.485 2.435 54.735 3.445 ;
  LAYER M1 ;
        RECT 54.485 0.335 54.735 1.345 ;
  LAYER M1 ;
        RECT 54.055 3.695 54.305 7.225 ;
  LAYER M1 ;
        RECT 54.915 3.695 55.165 7.225 ;
  LAYER M1 ;
        RECT 55.345 3.695 55.595 7.225 ;
  LAYER M1 ;
        RECT 55.345 2.435 55.595 3.445 ;
  LAYER M1 ;
        RECT 55.345 0.335 55.595 1.345 ;
  LAYER M1 ;
        RECT 55.775 3.695 56.025 7.225 ;
  LAYER M2 ;
        RECT 54.44 0.7 55.64 0.98 ;
  LAYER M2 ;
        RECT 54.01 6.58 56.07 6.86 ;
  LAYER M2 ;
        RECT 54.44 7 55.64 7.28 ;
  LAYER M2 ;
        RECT 54.44 2.8 55.64 3.08 ;
  LAYER M3 ;
        RECT 55.33 0.68 55.61 6.88 ;
  LAYER M1 ;
        RECT 39.005 7.895 39.255 11.425 ;
  LAYER M1 ;
        RECT 39.005 11.675 39.255 12.685 ;
  LAYER M1 ;
        RECT 39.005 13.775 39.255 14.785 ;
  LAYER M1 ;
        RECT 38.575 7.895 38.825 11.425 ;
  LAYER M1 ;
        RECT 39.435 7.895 39.685 11.425 ;
  LAYER M1 ;
        RECT 39.865 7.895 40.115 11.425 ;
  LAYER M1 ;
        RECT 39.865 11.675 40.115 12.685 ;
  LAYER M1 ;
        RECT 39.865 13.775 40.115 14.785 ;
  LAYER M1 ;
        RECT 40.295 7.895 40.545 11.425 ;
  LAYER M2 ;
        RECT 38.96 14.14 40.16 14.42 ;
  LAYER M2 ;
        RECT 38.53 8.26 40.59 8.54 ;
  LAYER M2 ;
        RECT 38.96 7.84 40.16 8.12 ;
  LAYER M2 ;
        RECT 38.96 12.04 40.16 12.32 ;
  LAYER M3 ;
        RECT 39.85 8.24 40.13 14.44 ;
  LAYER M1 ;
        RECT 39.865 3.695 40.115 7.225 ;
  LAYER M1 ;
        RECT 39.865 2.435 40.115 3.445 ;
  LAYER M1 ;
        RECT 39.865 0.335 40.115 1.345 ;
  LAYER M1 ;
        RECT 39.435 3.695 39.685 7.225 ;
  LAYER M1 ;
        RECT 40.295 3.695 40.545 7.225 ;
  LAYER M1 ;
        RECT 40.725 3.695 40.975 7.225 ;
  LAYER M1 ;
        RECT 40.725 2.435 40.975 3.445 ;
  LAYER M1 ;
        RECT 40.725 0.335 40.975 1.345 ;
  LAYER M1 ;
        RECT 41.155 3.695 41.405 7.225 ;
  LAYER M2 ;
        RECT 39.82 0.7 41.02 0.98 ;
  LAYER M2 ;
        RECT 39.82 7 41.02 7.28 ;
  LAYER M2 ;
        RECT 39.82 2.8 41.02 3.08 ;
  LAYER M2 ;
        RECT 39.39 6.58 41.45 6.86 ;
  LAYER M1 ;
        RECT 43.305 3.695 43.555 7.225 ;
  LAYER M1 ;
        RECT 43.305 2.435 43.555 3.445 ;
  LAYER M1 ;
        RECT 43.305 0.335 43.555 1.345 ;
  LAYER M1 ;
        RECT 42.875 3.695 43.125 7.225 ;
  LAYER M1 ;
        RECT 43.735 3.695 43.985 7.225 ;
  LAYER M1 ;
        RECT 44.165 3.695 44.415 7.225 ;
  LAYER M1 ;
        RECT 44.165 2.435 44.415 3.445 ;
  LAYER M1 ;
        RECT 44.165 0.335 44.415 1.345 ;
  LAYER M1 ;
        RECT 44.595 3.695 44.845 7.225 ;
  LAYER M2 ;
        RECT 43.26 0.7 44.46 0.98 ;
  LAYER M2 ;
        RECT 43.26 7 44.46 7.28 ;
  LAYER M2 ;
        RECT 43.26 2.8 44.46 3.08 ;
  LAYER M2 ;
        RECT 42.83 6.58 44.89 6.86 ;
  LAYER M2 ;
        RECT 24.34 7 25.54 7.28 ;
  LAYER M2 ;
        RECT 24.34 8.26 25.54 8.54 ;
  LAYER M2 ;
        RECT 28.64 2.8 29.84 3.08 ;
  LAYER M2 ;
        RECT 28.64 12.04 29.84 12.32 ;
  LAYER M2 ;
        RECT 29.08 2.8 29.4 3.08 ;
  LAYER M3 ;
        RECT 29.1 2.94 29.38 12.18 ;
  LAYER M2 ;
        RECT 29.08 12.04 29.4 12.32 ;
  LAYER M2 ;
        RECT 24.78 7 25.1 7.28 ;
  LAYER M3 ;
        RECT 24.8 7.14 25.08 8.4 ;
  LAYER M2 ;
        RECT 24.78 8.26 25.1 8.54 ;
  LAYER M3 ;
        RECT 24.8 7.375 25.08 7.745 ;
  LAYER M2 ;
        RECT 24.94 7.42 29.24 7.7 ;
  LAYER M3 ;
        RECT 29.1 7.375 29.38 7.745 ;
  LAYER M2 ;
        RECT 24.78 7 25.1 7.28 ;
  LAYER M3 ;
        RECT 24.8 6.98 25.08 7.3 ;
  LAYER M2 ;
        RECT 24.78 8.26 25.1 8.54 ;
  LAYER M3 ;
        RECT 24.8 8.24 25.08 8.56 ;
  LAYER M2 ;
        RECT 24.78 7 25.1 7.28 ;
  LAYER M3 ;
        RECT 24.8 6.98 25.08 7.3 ;
  LAYER M2 ;
        RECT 24.78 8.26 25.1 8.54 ;
  LAYER M3 ;
        RECT 24.8 8.24 25.08 8.56 ;
  LAYER M2 ;
        RECT 24.78 7 25.1 7.28 ;
  LAYER M3 ;
        RECT 24.8 6.98 25.08 7.3 ;
  LAYER M2 ;
        RECT 24.78 7.42 25.1 7.7 ;
  LAYER M3 ;
        RECT 24.8 7.4 25.08 7.72 ;
  LAYER M2 ;
        RECT 24.78 8.26 25.1 8.54 ;
  LAYER M3 ;
        RECT 24.8 8.24 25.08 8.56 ;
  LAYER M2 ;
        RECT 29.08 7.42 29.4 7.7 ;
  LAYER M3 ;
        RECT 29.1 7.4 29.38 7.72 ;
  LAYER M2 ;
        RECT 24.78 7 25.1 7.28 ;
  LAYER M3 ;
        RECT 24.8 6.98 25.08 7.3 ;
  LAYER M2 ;
        RECT 24.78 7.42 25.1 7.7 ;
  LAYER M3 ;
        RECT 24.8 7.4 25.08 7.72 ;
  LAYER M2 ;
        RECT 24.78 8.26 25.1 8.54 ;
  LAYER M3 ;
        RECT 24.8 8.24 25.08 8.56 ;
  LAYER M2 ;
        RECT 29.08 7.42 29.4 7.7 ;
  LAYER M3 ;
        RECT 29.1 7.4 29.38 7.72 ;
  LAYER M2 ;
        RECT 35.52 2.8 36.72 3.08 ;
  LAYER M2 ;
        RECT 35.52 12.04 36.72 12.32 ;
  LAYER M2 ;
        RECT 35.53 2.8 35.85 3.08 ;
  LAYER M3 ;
        RECT 35.55 2.94 35.83 12.18 ;
  LAYER M2 ;
        RECT 35.53 12.04 35.85 12.32 ;
  LAYER M2 ;
        RECT 32.08 7 33.28 7.28 ;
  LAYER M2 ;
        RECT 32.08 7.84 33.28 8.12 ;
  LAYER M2 ;
        RECT 32.52 7 32.84 7.28 ;
  LAYER M3 ;
        RECT 32.54 7.14 32.82 7.98 ;
  LAYER M2 ;
        RECT 32.52 7.84 32.84 8.12 ;
  LAYER M3 ;
        RECT 35.55 7.375 35.83 7.745 ;
  LAYER M2 ;
        RECT 32.68 7.42 35.69 7.7 ;
  LAYER M3 ;
        RECT 32.54 7.375 32.82 7.745 ;
  LAYER M2 ;
        RECT 32.52 7.42 32.84 7.7 ;
  LAYER M3 ;
        RECT 32.54 7.4 32.82 7.72 ;
  LAYER M2 ;
        RECT 35.53 7.42 35.85 7.7 ;
  LAYER M3 ;
        RECT 35.55 7.4 35.83 7.72 ;
  LAYER M2 ;
        RECT 32.52 7.42 32.84 7.7 ;
  LAYER M3 ;
        RECT 32.54 7.4 32.82 7.72 ;
  LAYER M2 ;
        RECT 35.53 7.42 35.85 7.7 ;
  LAYER M3 ;
        RECT 35.55 7.4 35.83 7.72 ;
  LAYER M2 ;
        RECT 20.9 7 22.1 7.28 ;
  LAYER M3 ;
        RECT 24.37 7.82 24.65 12.34 ;
  LAYER M2 ;
        RECT 21.93 7 23.65 7.28 ;
  LAYER M3 ;
        RECT 23.51 7.14 23.79 7.56 ;
  LAYER M4 ;
        RECT 23.65 7.16 24.51 7.96 ;
  LAYER M3 ;
        RECT 24.37 7.56 24.65 7.98 ;
  LAYER M2 ;
        RECT 23.49 7 23.81 7.28 ;
  LAYER M3 ;
        RECT 23.51 6.98 23.79 7.3 ;
  LAYER M3 ;
        RECT 23.51 7.375 23.79 7.745 ;
  LAYER M4 ;
        RECT 23.485 7.16 23.815 7.96 ;
  LAYER M3 ;
        RECT 24.37 7.375 24.65 7.745 ;
  LAYER M4 ;
        RECT 24.345 7.16 24.675 7.96 ;
  LAYER M2 ;
        RECT 23.49 7 23.81 7.28 ;
  LAYER M3 ;
        RECT 23.51 6.98 23.79 7.3 ;
  LAYER M3 ;
        RECT 23.51 7.375 23.79 7.745 ;
  LAYER M4 ;
        RECT 23.485 7.16 23.815 7.96 ;
  LAYER M3 ;
        RECT 24.37 7.375 24.65 7.745 ;
  LAYER M4 ;
        RECT 24.345 7.16 24.675 7.96 ;
  LAYER M2 ;
        RECT 20.47 6.58 22.53 6.86 ;
  LAYER M2 ;
        RECT 20.04 7.84 21.24 8.12 ;
  LAYER M2 ;
        RECT 23.91 6.58 25.97 6.86 ;
  LAYER M2 ;
        RECT 20.48 6.58 20.8 6.86 ;
  LAYER M3 ;
        RECT 20.5 6.72 20.78 7.98 ;
  LAYER M2 ;
        RECT 20.48 7.84 20.8 8.12 ;
  LAYER M2 ;
        RECT 22.36 6.58 24.08 6.86 ;
  LAYER M2 ;
        RECT 20.48 6.58 20.8 6.86 ;
  LAYER M3 ;
        RECT 20.5 6.56 20.78 6.88 ;
  LAYER M2 ;
        RECT 20.48 7.84 20.8 8.12 ;
  LAYER M3 ;
        RECT 20.5 7.82 20.78 8.14 ;
  LAYER M2 ;
        RECT 20.48 6.58 20.8 6.86 ;
  LAYER M3 ;
        RECT 20.5 6.56 20.78 6.88 ;
  LAYER M2 ;
        RECT 20.48 7.84 20.8 8.12 ;
  LAYER M3 ;
        RECT 20.5 7.82 20.78 8.14 ;
  LAYER M2 ;
        RECT 20.48 6.58 20.8 6.86 ;
  LAYER M3 ;
        RECT 20.5 6.56 20.78 6.88 ;
  LAYER M2 ;
        RECT 20.48 7.84 20.8 8.12 ;
  LAYER M3 ;
        RECT 20.5 7.82 20.78 8.14 ;
  LAYER M2 ;
        RECT 20.48 6.58 20.8 6.86 ;
  LAYER M3 ;
        RECT 20.5 6.56 20.78 6.88 ;
  LAYER M2 ;
        RECT 20.48 7.84 20.8 8.12 ;
  LAYER M3 ;
        RECT 20.5 7.82 20.78 8.14 ;
  LAYER M2 ;
        RECT 32.08 2.8 33.28 3.08 ;
  LAYER M2 ;
        RECT 28.64 7 29.84 7.28 ;
  LAYER M2 ;
        RECT 28.64 7.84 29.84 8.12 ;
  LAYER M2 ;
        RECT 32.08 12.04 33.28 12.32 ;
  LAYER M2 ;
        RECT 30.96 2.8 32.25 3.08 ;
  LAYER M1 ;
        RECT 30.835 2.94 31.085 7.14 ;
  LAYER M2 ;
        RECT 29.67 7 30.96 7.28 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 7.14 29.81 7.98 ;
  LAYER M2 ;
        RECT 29.51 7.84 29.83 8.12 ;
  LAYER M1 ;
        RECT 30.835 7.14 31.085 12.18 ;
  LAYER M2 ;
        RECT 30.96 12.04 32.25 12.32 ;
  LAYER M1 ;
        RECT 30.835 2.855 31.085 3.025 ;
  LAYER M2 ;
        RECT 30.79 2.8 31.13 3.08 ;
  LAYER M1 ;
        RECT 30.835 7.055 31.085 7.225 ;
  LAYER M2 ;
        RECT 30.79 7 31.13 7.28 ;
  LAYER M1 ;
        RECT 30.835 2.855 31.085 3.025 ;
  LAYER M2 ;
        RECT 30.79 2.8 31.13 3.08 ;
  LAYER M1 ;
        RECT 30.835 7.055 31.085 7.225 ;
  LAYER M2 ;
        RECT 30.79 7 31.13 7.28 ;
  LAYER M1 ;
        RECT 30.835 2.855 31.085 3.025 ;
  LAYER M2 ;
        RECT 30.79 2.8 31.13 3.08 ;
  LAYER M1 ;
        RECT 30.835 7.055 31.085 7.225 ;
  LAYER M2 ;
        RECT 30.79 7 31.13 7.28 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 6.98 29.81 7.3 ;
  LAYER M2 ;
        RECT 29.51 7.84 29.83 8.12 ;
  LAYER M3 ;
        RECT 29.53 7.82 29.81 8.14 ;
  LAYER M1 ;
        RECT 30.835 2.855 31.085 3.025 ;
  LAYER M2 ;
        RECT 30.79 2.8 31.13 3.08 ;
  LAYER M1 ;
        RECT 30.835 7.055 31.085 7.225 ;
  LAYER M2 ;
        RECT 30.79 7 31.13 7.28 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 6.98 29.81 7.3 ;
  LAYER M2 ;
        RECT 29.51 7.84 29.83 8.12 ;
  LAYER M3 ;
        RECT 29.53 7.82 29.81 8.14 ;
  LAYER M1 ;
        RECT 30.835 2.855 31.085 3.025 ;
  LAYER M2 ;
        RECT 30.79 2.8 31.13 3.08 ;
  LAYER M1 ;
        RECT 30.835 7.055 31.085 7.225 ;
  LAYER M2 ;
        RECT 30.79 7 31.13 7.28 ;
  LAYER M1 ;
        RECT 30.835 12.095 31.085 12.265 ;
  LAYER M2 ;
        RECT 30.79 12.04 31.13 12.32 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 6.98 29.81 7.3 ;
  LAYER M2 ;
        RECT 29.51 7.84 29.83 8.12 ;
  LAYER M3 ;
        RECT 29.53 7.82 29.81 8.14 ;
  LAYER M1 ;
        RECT 30.835 2.855 31.085 3.025 ;
  LAYER M2 ;
        RECT 30.79 2.8 31.13 3.08 ;
  LAYER M1 ;
        RECT 30.835 7.055 31.085 7.225 ;
  LAYER M2 ;
        RECT 30.79 7 31.13 7.28 ;
  LAYER M1 ;
        RECT 30.835 12.095 31.085 12.265 ;
  LAYER M2 ;
        RECT 30.79 12.04 31.13 12.32 ;
  LAYER M2 ;
        RECT 29.51 7 29.83 7.28 ;
  LAYER M3 ;
        RECT 29.53 6.98 29.81 7.3 ;
  LAYER M2 ;
        RECT 29.51 7.84 29.83 8.12 ;
  LAYER M3 ;
        RECT 29.53 7.82 29.81 8.14 ;
  LAYER M1 ;
        RECT 29.545 7.895 29.795 11.425 ;
  LAYER M1 ;
        RECT 29.545 11.675 29.795 12.685 ;
  LAYER M1 ;
        RECT 29.545 13.775 29.795 14.785 ;
  LAYER M1 ;
        RECT 29.975 7.895 30.225 11.425 ;
  LAYER M1 ;
        RECT 29.115 7.895 29.365 11.425 ;
  LAYER M1 ;
        RECT 28.685 7.895 28.935 11.425 ;
  LAYER M1 ;
        RECT 28.685 11.675 28.935 12.685 ;
  LAYER M1 ;
        RECT 28.685 13.775 28.935 14.785 ;
  LAYER M1 ;
        RECT 28.255 7.895 28.505 11.425 ;
  LAYER M2 ;
        RECT 28.64 14.14 29.84 14.42 ;
  LAYER M2 ;
        RECT 28.21 8.26 30.27 8.54 ;
  LAYER M2 ;
        RECT 28.64 7.84 29.84 8.12 ;
  LAYER M2 ;
        RECT 28.64 12.04 29.84 12.32 ;
  LAYER M3 ;
        RECT 28.67 8.24 28.95 14.44 ;
  LAYER M1 ;
        RECT 32.985 7.895 33.235 11.425 ;
  LAYER M1 ;
        RECT 32.985 11.675 33.235 12.685 ;
  LAYER M1 ;
        RECT 32.985 13.775 33.235 14.785 ;
  LAYER M1 ;
        RECT 33.415 7.895 33.665 11.425 ;
  LAYER M1 ;
        RECT 32.555 7.895 32.805 11.425 ;
  LAYER M1 ;
        RECT 32.125 7.895 32.375 11.425 ;
  LAYER M1 ;
        RECT 32.125 11.675 32.375 12.685 ;
  LAYER M1 ;
        RECT 32.125 13.775 32.375 14.785 ;
  LAYER M1 ;
        RECT 31.695 7.895 31.945 11.425 ;
  LAYER M2 ;
        RECT 32.08 14.14 33.28 14.42 ;
  LAYER M2 ;
        RECT 31.65 8.26 33.71 8.54 ;
  LAYER M2 ;
        RECT 32.08 7.84 33.28 8.12 ;
  LAYER M2 ;
        RECT 32.08 12.04 33.28 12.32 ;
  LAYER M3 ;
        RECT 32.11 8.24 32.39 14.44 ;
  LAYER M1 ;
        RECT 29.545 3.695 29.795 7.225 ;
  LAYER M1 ;
        RECT 29.545 2.435 29.795 3.445 ;
  LAYER M1 ;
        RECT 29.545 0.335 29.795 1.345 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M1 ;
        RECT 29.115 3.695 29.365 7.225 ;
  LAYER M1 ;
        RECT 28.685 3.695 28.935 7.225 ;
  LAYER M1 ;
        RECT 28.685 2.435 28.935 3.445 ;
  LAYER M1 ;
        RECT 28.685 0.335 28.935 1.345 ;
  LAYER M1 ;
        RECT 28.255 3.695 28.505 7.225 ;
  LAYER M2 ;
        RECT 28.64 0.7 29.84 0.98 ;
  LAYER M2 ;
        RECT 28.21 6.58 30.27 6.86 ;
  LAYER M2 ;
        RECT 28.64 7 29.84 7.28 ;
  LAYER M2 ;
        RECT 28.64 2.8 29.84 3.08 ;
  LAYER M3 ;
        RECT 28.67 0.68 28.95 6.88 ;
  LAYER M1 ;
        RECT 32.985 3.695 33.235 7.225 ;
  LAYER M1 ;
        RECT 32.985 2.435 33.235 3.445 ;
  LAYER M1 ;
        RECT 32.985 0.335 33.235 1.345 ;
  LAYER M1 ;
        RECT 33.415 3.695 33.665 7.225 ;
  LAYER M1 ;
        RECT 32.555 3.695 32.805 7.225 ;
  LAYER M1 ;
        RECT 32.125 3.695 32.375 7.225 ;
  LAYER M1 ;
        RECT 32.125 2.435 32.375 3.445 ;
  LAYER M1 ;
        RECT 32.125 0.335 32.375 1.345 ;
  LAYER M1 ;
        RECT 31.695 3.695 31.945 7.225 ;
  LAYER M2 ;
        RECT 32.08 0.7 33.28 0.98 ;
  LAYER M2 ;
        RECT 31.65 6.58 33.71 6.86 ;
  LAYER M2 ;
        RECT 32.08 7 33.28 7.28 ;
  LAYER M2 ;
        RECT 32.08 2.8 33.28 3.08 ;
  LAYER M3 ;
        RECT 32.11 0.68 32.39 6.88 ;
  LAYER M1 ;
        RECT 23.525 7.895 23.775 11.425 ;
  LAYER M1 ;
        RECT 23.525 11.675 23.775 12.685 ;
  LAYER M1 ;
        RECT 23.525 13.775 23.775 14.785 ;
  LAYER M1 ;
        RECT 23.095 7.895 23.345 11.425 ;
  LAYER M1 ;
        RECT 23.955 7.895 24.205 11.425 ;
  LAYER M1 ;
        RECT 24.385 7.895 24.635 11.425 ;
  LAYER M1 ;
        RECT 24.385 11.675 24.635 12.685 ;
  LAYER M1 ;
        RECT 24.385 13.775 24.635 14.785 ;
  LAYER M1 ;
        RECT 24.815 7.895 25.065 11.425 ;
  LAYER M1 ;
        RECT 25.245 7.895 25.495 11.425 ;
  LAYER M1 ;
        RECT 25.245 11.675 25.495 12.685 ;
  LAYER M1 ;
        RECT 25.245 13.775 25.495 14.785 ;
  LAYER M1 ;
        RECT 25.675 7.895 25.925 11.425 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 11.425 ;
  LAYER M1 ;
        RECT 26.105 11.675 26.355 12.685 ;
  LAYER M1 ;
        RECT 26.105 13.775 26.355 14.785 ;
  LAYER M1 ;
        RECT 26.535 7.895 26.785 11.425 ;
  LAYER M2 ;
        RECT 23.48 12.04 26.4 12.32 ;
  LAYER M2 ;
        RECT 23.48 7.84 26.4 8.12 ;
  LAYER M2 ;
        RECT 23.48 14.14 26.4 14.42 ;
  LAYER M2 ;
        RECT 23.05 8.68 26.83 8.96 ;
  LAYER M3 ;
        RECT 24.37 7.82 24.65 12.34 ;
  LAYER M2 ;
        RECT 24.34 8.26 25.54 8.54 ;
  LAYER M3 ;
        RECT 25.23 8.66 25.51 14.44 ;
  LAYER M1 ;
        RECT 35.565 7.895 35.815 11.425 ;
  LAYER M1 ;
        RECT 35.565 11.675 35.815 12.685 ;
  LAYER M1 ;
        RECT 35.565 13.775 35.815 14.785 ;
  LAYER M1 ;
        RECT 35.135 7.895 35.385 11.425 ;
  LAYER M1 ;
        RECT 35.995 7.895 36.245 11.425 ;
  LAYER M1 ;
        RECT 36.425 7.895 36.675 11.425 ;
  LAYER M1 ;
        RECT 36.425 11.675 36.675 12.685 ;
  LAYER M1 ;
        RECT 36.425 13.775 36.675 14.785 ;
  LAYER M1 ;
        RECT 36.855 7.895 37.105 11.425 ;
  LAYER M2 ;
        RECT 35.52 14.14 36.72 14.42 ;
  LAYER M2 ;
        RECT 35.09 8.26 37.15 8.54 ;
  LAYER M2 ;
        RECT 35.52 7.84 36.72 8.12 ;
  LAYER M2 ;
        RECT 35.52 12.04 36.72 12.32 ;
  LAYER M3 ;
        RECT 36.41 8.24 36.69 14.44 ;
  LAYER M1 ;
        RECT 35.565 3.695 35.815 7.225 ;
  LAYER M1 ;
        RECT 35.565 2.435 35.815 3.445 ;
  LAYER M1 ;
        RECT 35.565 0.335 35.815 1.345 ;
  LAYER M1 ;
        RECT 35.135 3.695 35.385 7.225 ;
  LAYER M1 ;
        RECT 35.995 3.695 36.245 7.225 ;
  LAYER M1 ;
        RECT 36.425 3.695 36.675 7.225 ;
  LAYER M1 ;
        RECT 36.425 2.435 36.675 3.445 ;
  LAYER M1 ;
        RECT 36.425 0.335 36.675 1.345 ;
  LAYER M1 ;
        RECT 36.855 3.695 37.105 7.225 ;
  LAYER M2 ;
        RECT 35.52 0.7 36.72 0.98 ;
  LAYER M2 ;
        RECT 35.09 6.58 37.15 6.86 ;
  LAYER M2 ;
        RECT 35.52 7 36.72 7.28 ;
  LAYER M2 ;
        RECT 35.52 2.8 36.72 3.08 ;
  LAYER M3 ;
        RECT 36.41 0.68 36.69 6.88 ;
  LAYER M1 ;
        RECT 20.085 7.895 20.335 11.425 ;
  LAYER M1 ;
        RECT 20.085 11.675 20.335 12.685 ;
  LAYER M1 ;
        RECT 20.085 13.775 20.335 14.785 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M1 ;
        RECT 20.515 7.895 20.765 11.425 ;
  LAYER M1 ;
        RECT 20.945 7.895 21.195 11.425 ;
  LAYER M1 ;
        RECT 20.945 11.675 21.195 12.685 ;
  LAYER M1 ;
        RECT 20.945 13.775 21.195 14.785 ;
  LAYER M1 ;
        RECT 21.375 7.895 21.625 11.425 ;
  LAYER M2 ;
        RECT 20.04 14.14 21.24 14.42 ;
  LAYER M2 ;
        RECT 19.61 8.26 21.67 8.54 ;
  LAYER M2 ;
        RECT 20.04 7.84 21.24 8.12 ;
  LAYER M2 ;
        RECT 20.04 12.04 21.24 12.32 ;
  LAYER M3 ;
        RECT 20.93 8.24 21.21 14.44 ;
  LAYER M1 ;
        RECT 20.945 3.695 21.195 7.225 ;
  LAYER M1 ;
        RECT 20.945 2.435 21.195 3.445 ;
  LAYER M1 ;
        RECT 20.945 0.335 21.195 1.345 ;
  LAYER M1 ;
        RECT 20.515 3.695 20.765 7.225 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M1 ;
        RECT 21.805 3.695 22.055 7.225 ;
  LAYER M1 ;
        RECT 21.805 2.435 22.055 3.445 ;
  LAYER M1 ;
        RECT 21.805 0.335 22.055 1.345 ;
  LAYER M1 ;
        RECT 22.235 3.695 22.485 7.225 ;
  LAYER M2 ;
        RECT 20.9 0.7 22.1 0.98 ;
  LAYER M2 ;
        RECT 20.9 7 22.1 7.28 ;
  LAYER M2 ;
        RECT 20.9 2.8 22.1 3.08 ;
  LAYER M2 ;
        RECT 20.47 6.58 22.53 6.86 ;
  LAYER M1 ;
        RECT 24.385 3.695 24.635 7.225 ;
  LAYER M1 ;
        RECT 24.385 2.435 24.635 3.445 ;
  LAYER M1 ;
        RECT 24.385 0.335 24.635 1.345 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M2 ;
        RECT 24.34 0.7 25.54 0.98 ;
  LAYER M2 ;
        RECT 24.34 7 25.54 7.28 ;
  LAYER M2 ;
        RECT 24.34 2.8 25.54 3.08 ;
  LAYER M2 ;
        RECT 23.91 6.58 25.97 6.86 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M2 ;
        RECT 8.44 2.8 8.76 3.08 ;
  LAYER M3 ;
        RECT 8.46 2.94 8.74 12.18 ;
  LAYER M2 ;
        RECT 8.44 12.04 8.76 12.32 ;
  LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 12.3 8.26 13.5 8.54 ;
  LAYER M3 ;
        RECT 8.46 7.375 8.74 7.745 ;
  LAYER M2 ;
        RECT 8.6 7.42 9.89 7.7 ;
  LAYER M1 ;
        RECT 9.765 7.14 10.015 7.56 ;
  LAYER M2 ;
        RECT 9.89 7 12.47 7.28 ;
  LAYER M2 ;
        RECT 12.74 7 13.06 7.28 ;
  LAYER M3 ;
        RECT 12.76 7.14 13.04 8.4 ;
  LAYER M2 ;
        RECT 12.74 8.26 13.06 8.54 ;
  LAYER M1 ;
        RECT 9.765 7.055 10.015 7.225 ;
  LAYER M2 ;
        RECT 9.72 7 10.06 7.28 ;
  LAYER M1 ;
        RECT 9.765 7.475 10.015 7.645 ;
  LAYER M2 ;
        RECT 9.72 7.42 10.06 7.7 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M1 ;
        RECT 9.765 7.055 10.015 7.225 ;
  LAYER M2 ;
        RECT 9.72 7 10.06 7.28 ;
  LAYER M1 ;
        RECT 9.765 7.475 10.015 7.645 ;
  LAYER M2 ;
        RECT 9.72 7.42 10.06 7.7 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M1 ;
        RECT 9.765 7.055 10.015 7.225 ;
  LAYER M2 ;
        RECT 9.72 7 10.06 7.28 ;
  LAYER M1 ;
        RECT 9.765 7.475 10.015 7.645 ;
  LAYER M2 ;
        RECT 9.72 7.42 10.06 7.7 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 12.74 7 13.06 7.28 ;
  LAYER M3 ;
        RECT 12.76 6.98 13.04 7.3 ;
  LAYER M2 ;
        RECT 12.74 8.26 13.06 8.54 ;
  LAYER M3 ;
        RECT 12.76 8.24 13.04 8.56 ;
  LAYER M1 ;
        RECT 9.765 7.055 10.015 7.225 ;
  LAYER M2 ;
        RECT 9.72 7 10.06 7.28 ;
  LAYER M1 ;
        RECT 9.765 7.475 10.015 7.645 ;
  LAYER M2 ;
        RECT 9.72 7.42 10.06 7.7 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 12.74 7 13.06 7.28 ;
  LAYER M3 ;
        RECT 12.76 6.98 13.04 7.3 ;
  LAYER M2 ;
        RECT 12.74 8.26 13.06 8.54 ;
  LAYER M3 ;
        RECT 12.76 8.24 13.04 8.56 ;
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 1.99 2.8 2.31 3.08 ;
  LAYER M3 ;
        RECT 2.01 2.94 2.29 12.18 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M2 ;
        RECT 4.56 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 4.56 7.84 5.76 8.12 ;
  LAYER M2 ;
        RECT 5 7 5.32 7.28 ;
  LAYER M3 ;
        RECT 5.02 7.14 5.3 7.98 ;
  LAYER M2 ;
        RECT 5 7.84 5.32 8.12 ;
  LAYER M3 ;
        RECT 2.01 7.375 2.29 7.745 ;
  LAYER M2 ;
        RECT 2.15 7.42 5.16 7.7 ;
  LAYER M3 ;
        RECT 5.02 7.375 5.3 7.745 ;
  LAYER M2 ;
        RECT 1.99 7.42 2.31 7.7 ;
  LAYER M3 ;
        RECT 2.01 7.4 2.29 7.72 ;
  LAYER M2 ;
        RECT 5 7.42 5.32 7.7 ;
  LAYER M3 ;
        RECT 5.02 7.4 5.3 7.72 ;
  LAYER M2 ;
        RECT 1.99 7.42 2.31 7.7 ;
  LAYER M3 ;
        RECT 2.01 7.4 2.29 7.72 ;
  LAYER M2 ;
        RECT 5 7.42 5.32 7.7 ;
  LAYER M3 ;
        RECT 5.02 7.4 5.3 7.72 ;
  LAYER M3 ;
        RECT 13.19 7.82 13.47 12.34 ;
  LAYER M2 ;
        RECT 15.74 7 16.94 7.28 ;
  LAYER M3 ;
        RECT 13.19 7.56 13.47 7.98 ;
  LAYER M2 ;
        RECT 13.33 7.42 15.05 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.14 15.175 7.56 ;
  LAYER M2 ;
        RECT 15.05 7 15.91 7.28 ;
  LAYER M1 ;
        RECT 14.925 7.055 15.175 7.225 ;
  LAYER M2 ;
        RECT 14.88 7 15.22 7.28 ;
  LAYER M1 ;
        RECT 14.925 7.475 15.175 7.645 ;
  LAYER M2 ;
        RECT 14.88 7.42 15.22 7.7 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M1 ;
        RECT 14.925 7.055 15.175 7.225 ;
  LAYER M2 ;
        RECT 14.88 7 15.22 7.28 ;
  LAYER M1 ;
        RECT 14.925 7.475 15.175 7.645 ;
  LAYER M2 ;
        RECT 14.88 7.42 15.22 7.7 ;
  LAYER M2 ;
        RECT 13.17 7.42 13.49 7.7 ;
  LAYER M3 ;
        RECT 13.19 7.4 13.47 7.72 ;
  LAYER M2 ;
        RECT 11.87 6.58 13.93 6.86 ;
  LAYER M2 ;
        RECT 15.31 6.58 17.37 6.86 ;
  LAYER M2 ;
        RECT 16.6 7.84 17.8 8.12 ;
  LAYER M2 ;
        RECT 13.76 6.58 15.48 6.86 ;
  LAYER M2 ;
        RECT 17.04 6.58 17.36 6.86 ;
  LAYER M3 ;
        RECT 17.06 6.72 17.34 7.98 ;
  LAYER M2 ;
        RECT 17.04 7.84 17.36 8.12 ;
  LAYER M2 ;
        RECT 17.04 6.58 17.36 6.86 ;
  LAYER M3 ;
        RECT 17.06 6.56 17.34 6.88 ;
  LAYER M2 ;
        RECT 17.04 7.84 17.36 8.12 ;
  LAYER M3 ;
        RECT 17.06 7.82 17.34 8.14 ;
  LAYER M2 ;
        RECT 17.04 6.58 17.36 6.86 ;
  LAYER M3 ;
        RECT 17.06 6.56 17.34 6.88 ;
  LAYER M2 ;
        RECT 17.04 7.84 17.36 8.12 ;
  LAYER M3 ;
        RECT 17.06 7.82 17.34 8.14 ;
  LAYER M2 ;
        RECT 4.56 2.8 5.76 3.08 ;
  LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 4.56 12.04 5.76 12.32 ;
  LAYER M2 ;
        RECT 5.59 2.8 6.88 3.08 ;
  LAYER M1 ;
        RECT 6.755 2.94 7.005 7.14 ;
  LAYER M2 ;
        RECT 6.88 7 8.17 7.28 ;
  LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
  LAYER M3 ;
        RECT 8.03 7.14 8.31 7.98 ;
  LAYER M2 ;
        RECT 8.01 7.84 8.33 8.12 ;
  LAYER M1 ;
        RECT 6.755 7.14 7.005 12.18 ;
  LAYER M2 ;
        RECT 5.59 12.04 6.88 12.32 ;
  LAYER M1 ;
        RECT 6.755 2.855 7.005 3.025 ;
  LAYER M2 ;
        RECT 6.71 2.8 7.05 3.08 ;
  LAYER M1 ;
        RECT 6.755 7.055 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 7 7.05 7.28 ;
  LAYER M1 ;
        RECT 6.755 2.855 7.005 3.025 ;
  LAYER M2 ;
        RECT 6.71 2.8 7.05 3.08 ;
  LAYER M1 ;
        RECT 6.755 7.055 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 7 7.05 7.28 ;
  LAYER M1 ;
        RECT 6.755 2.855 7.005 3.025 ;
  LAYER M2 ;
        RECT 6.71 2.8 7.05 3.08 ;
  LAYER M1 ;
        RECT 6.755 7.055 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 7 7.05 7.28 ;
  LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
  LAYER M3 ;
        RECT 8.03 6.98 8.31 7.3 ;
  LAYER M2 ;
        RECT 8.01 7.84 8.33 8.12 ;
  LAYER M3 ;
        RECT 8.03 7.82 8.31 8.14 ;
  LAYER M1 ;
        RECT 6.755 2.855 7.005 3.025 ;
  LAYER M2 ;
        RECT 6.71 2.8 7.05 3.08 ;
  LAYER M1 ;
        RECT 6.755 7.055 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 7 7.05 7.28 ;
  LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
  LAYER M3 ;
        RECT 8.03 6.98 8.31 7.3 ;
  LAYER M2 ;
        RECT 8.01 7.84 8.33 8.12 ;
  LAYER M3 ;
        RECT 8.03 7.82 8.31 8.14 ;
  LAYER M1 ;
        RECT 6.755 2.855 7.005 3.025 ;
  LAYER M2 ;
        RECT 6.71 2.8 7.05 3.08 ;
  LAYER M1 ;
        RECT 6.755 7.055 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 7 7.05 7.28 ;
  LAYER M1 ;
        RECT 6.755 12.095 7.005 12.265 ;
  LAYER M2 ;
        RECT 6.71 12.04 7.05 12.32 ;
  LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
  LAYER M3 ;
        RECT 8.03 6.98 8.31 7.3 ;
  LAYER M2 ;
        RECT 8.01 7.84 8.33 8.12 ;
  LAYER M3 ;
        RECT 8.03 7.82 8.31 8.14 ;
  LAYER M1 ;
        RECT 6.755 2.855 7.005 3.025 ;
  LAYER M2 ;
        RECT 6.71 2.8 7.05 3.08 ;
  LAYER M1 ;
        RECT 6.755 7.055 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 7 7.05 7.28 ;
  LAYER M1 ;
        RECT 6.755 12.095 7.005 12.265 ;
  LAYER M2 ;
        RECT 6.71 12.04 7.05 12.32 ;
  LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
  LAYER M3 ;
        RECT 8.03 6.98 8.31 7.3 ;
  LAYER M2 ;
        RECT 8.01 7.84 8.33 8.12 ;
  LAYER M3 ;
        RECT 8.03 7.82 8.31 8.14 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 14.785 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M2 ;
        RECT 8 14.14 9.2 14.42 ;
  LAYER M2 ;
        RECT 7.57 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M3 ;
        RECT 8.89 8.24 9.17 14.44 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 11.425 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 12.685 ;
  LAYER M1 ;
        RECT 4.605 13.775 4.855 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 11.425 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 11.425 ;
  LAYER M1 ;
        RECT 5.465 11.675 5.715 12.685 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M2 ;
        RECT 4.56 14.14 5.76 14.42 ;
  LAYER M2 ;
        RECT 4.13 8.26 6.19 8.54 ;
  LAYER M2 ;
        RECT 4.56 7.84 5.76 8.12 ;
  LAYER M2 ;
        RECT 4.56 12.04 5.76 12.32 ;
  LAYER M3 ;
        RECT 5.45 8.24 5.73 14.44 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 8 0.7 9.2 0.98 ;
  LAYER M2 ;
        RECT 7.57 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M3 ;
        RECT 8.89 0.68 9.17 6.88 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M2 ;
        RECT 4.56 0.7 5.76 0.98 ;
  LAYER M2 ;
        RECT 4.13 6.58 6.19 6.86 ;
  LAYER M2 ;
        RECT 4.56 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 4.56 2.8 5.76 3.08 ;
  LAYER M3 ;
        RECT 5.45 0.68 5.73 6.88 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 11.425 ;
  LAYER M1 ;
        RECT 13.205 11.675 13.455 12.685 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 14.785 ;
  LAYER M1 ;
        RECT 12.775 7.895 13.025 11.425 ;
  LAYER M1 ;
        RECT 12.345 7.895 12.595 11.425 ;
  LAYER M1 ;
        RECT 12.345 11.675 12.595 12.685 ;
  LAYER M1 ;
        RECT 12.345 13.775 12.595 14.785 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M2 ;
        RECT 11.44 12.04 14.36 12.32 ;
  LAYER M2 ;
        RECT 11.44 7.84 14.36 8.12 ;
  LAYER M2 ;
        RECT 11.44 14.14 14.36 14.42 ;
  LAYER M2 ;
        RECT 11.01 8.68 14.79 8.96 ;
  LAYER M3 ;
        RECT 13.19 7.82 13.47 12.34 ;
  LAYER M2 ;
        RECT 12.3 8.26 13.5 8.54 ;
  LAYER M3 ;
        RECT 12.33 8.66 12.61 14.44 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M2 ;
        RECT 1.12 14.14 2.32 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 2.75 8.54 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M3 ;
        RECT 1.15 8.24 1.43 14.44 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M2 ;
        RECT 1.12 0.7 2.32 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 2.75 6.86 ;
  LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M3 ;
        RECT 1.15 0.68 1.43 6.88 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 11.425 ;
  LAYER M1 ;
        RECT 17.505 11.675 17.755 12.685 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 14.785 ;
  LAYER M1 ;
        RECT 17.935 7.895 18.185 11.425 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 12.685 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 14.785 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M2 ;
        RECT 16.6 14.14 17.8 14.42 ;
  LAYER M2 ;
        RECT 16.17 8.26 18.23 8.54 ;
  LAYER M2 ;
        RECT 16.6 7.84 17.8 8.12 ;
  LAYER M2 ;
        RECT 16.6 12.04 17.8 12.32 ;
  LAYER M3 ;
        RECT 16.63 8.24 16.91 14.44 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M2 ;
        RECT 15.74 0.7 16.94 0.98 ;
  LAYER M2 ;
        RECT 15.74 7 16.94 7.28 ;
  LAYER M2 ;
        RECT 15.74 2.8 16.94 3.08 ;
  LAYER M2 ;
        RECT 15.31 6.58 17.37 6.86 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M2 ;
        RECT 12.3 0.7 13.5 0.98 ;
  LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
  LAYER M2 ;
        RECT 11.87 6.58 13.93 6.86 ;
  END 
END TWOBIT_FLASH_ADC
