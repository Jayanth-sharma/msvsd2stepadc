.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice  tt
X0 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=9e+11p pd=4.9e+06u as=9e+11p ps=4.9e+06u w=2e+06u l=150000u
X1 Vout Vin gnd gnd sky130_fd_pr__nfet_01v8 ad=4.5e+11p pd=2.9e+06u as=4.5e+11p ps=2.9e+06u w=1e+06u l=150000u


Vin Vin GND pulse(0 1.8 1n 1n 1n 4n 8n)
V2 Vdd GND 1.8


.tran 0.01n 60n
.control
run
.endc
.end

