magic
tech sky130A
magscale 1 2
timestamp 1677855779
<< locali >>
rect 61 2419 69 2453
rect 103 2419 111 2453
rect 61 605 111 2419
rect 61 571 69 605
rect 103 571 111 605
<< viali >>
rect 69 2419 103 2453
rect 69 571 103 605
<< metal1 >>
rect 52 2453 120 2464
rect 52 2419 69 2453
rect 103 2419 120 2453
rect 52 2408 120 2419
rect 140 1622 204 1624
rect 140 1570 146 1622
rect 198 1570 204 1622
rect 140 1568 204 1570
rect 140 1454 204 1456
rect 140 1402 146 1454
rect 198 1402 204 1454
rect 140 1400 204 1402
rect 52 605 120 616
rect 52 571 69 605
rect 103 571 120 605
rect 52 560 120 571
<< via1 >>
rect 146 1570 198 1622
rect 146 1402 198 1454
<< metal2 >>
rect 144 1622 200 1628
rect 144 1570 146 1622
rect 198 1570 200 1622
rect 144 1454 200 1570
rect 144 1402 146 1454
rect 198 1402 200 1454
rect 144 1396 200 1402
use NMOS_S_81537667_X1_Y1_1677853260_1677853264  NMOS_S_81537667_X1_Y1_1677853260_1677853264_0
timestamp 1677855779
transform 1 0 0 0 -1 1512
box 52 56 395 1482
use PMOS_4T_68898473_X1_Y1_1677853261_1677853264  PMOS_4T_68898473_X1_Y1_1677853261_1677853264_0
timestamp 1677855779
transform 1 0 0 0 1 1512
box 0 0 516 1512
<< end >>
