* SPICE3 file created from COMPARATOR_0.ext - technology: sky130A
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.subckt comparator VDD VSS VBIAS VIN VREF OUT
X0 VSS STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_2720_1484# VSS sky130_fd_pr__nfet_01v8 ad=2.7216e+12p pd=2.664e+07u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X1 m1_2720_1484# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 VSS STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_2720_1484# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 m1_2720_1484# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 VSS m1_1172_1316# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X5 STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_1172_1316# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 VSS m1_1172_1316# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_1172_1316# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 m1_2720_1484# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=3.192e+12p ps=3.112e+07u w=840000u l=150000u
X9 VDD STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_2720_1484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 m1_2720_1484# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 VDD STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_2720_1484# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_1172_1316# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X13 VDD m1_1172_1316# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_1172_1316# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 VDD m1_1172_1316# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 m1_688_1652# VREF m1_1172_1316# VSS sky130_fd_pr__nfet_01v8 ad=1.8312e+12p pd=1.78e+07u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X17 m1_1172_1316# VREF m1_688_1652# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18 m1_688_1652# VREF m1_1172_1316# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 m1_1172_1316# VREF m1_688_1652# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 m1_688_1652# NMOS_4T_77406006_X2_Y1_1679758483_1/a_200_252# m1_602_1568# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X21 m1_602_1568# NMOS_4T_77406006_X2_Y1_1679758483_1/a_200_252# m1_688_1652# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 m1_688_1652# NMOS_4T_77406006_X2_Y1_1679758483_1/a_200_252# m1_602_1568# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 m1_602_1568# NMOS_4T_77406006_X2_Y1_1679758483_1/a_200_252# m1_688_1652# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24 VDD m1_602_1568# m1_602_1568# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X25 m1_1172_1316# m1_602_1568# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X26 m1_602_1568# m1_602_1568# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 VDD m1_602_1568# m1_602_1568# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 VDD m1_602_1568# m1_1172_1316# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X29 m1_1172_1316# m1_602_1568# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X30 m1_602_1568# m1_602_1568# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 VDD m1_602_1568# m1_1172_1316# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X32 INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# m1_2720_1484# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X33 VDD m1_2720_1484# INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X34 INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# m1_2720_1484# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X35 VDD m1_2720_1484# INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X36 VSS m1_2720_1484# INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X37 INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# m1_2720_1484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X38 VSS m1_2720_1484# INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X39 INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# m1_2720_1484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X40 VSS NMOS_S_74334133_X2_Y1_1679758484_0/a_200_252# m1_688_1652# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X41 m1_688_1652# NMOS_S_74334133_X2_Y1_1679758484_0/a_200_252# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X42 VSS NMOS_S_74334133_X2_Y1_1679758484_0/a_200_252# m1_688_1652# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X43 m1_688_1652# NMOS_S_74334133_X2_Y1_1679758484_0/a_200_252# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 VREF VDD 0.03fF
C1 VREF m1_602_1568# 0.00fF
C2 VDD m1_2720_1484# 3.93fF
C3 VREF STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# 0.00fF
C4 VBIAS VDD 0.08fF
C5 m1_2720_1484# m1_602_1568# 0.00fF
C6 VBIAS m1_602_1568# 0.04fF
C7 m1_2720_1484# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# 0.57fF
C8 VREF m1_1172_1316# 0.26fF
C9 VDD m1_688_1652# 0.17fF
C10 m1_688_1652# m1_602_1568# 1.74fF
C11 m1_1172_1316# m1_2720_1484# 0.01fF
C12 m1_688_1652# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# 0.00fF
C13 VBIAS m1_1172_1316# 0.00fF
C14 m1_1172_1316# m1_688_1652# 1.38fF
C15 NMOS_4T_77406006_X2_Y1_1679758483_1/a_200_252# m1_602_1568# 0.22fF
C16 VDD OUT 0.15fF
C17 VREF m1_2720_1484# 0.00fF
C18 STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# OUT 0.00fF
C19 VIN VDD 0.00fF
C20 m1_1172_1316# OUT 0.00fF
C21 VIN m1_602_1568# 0.00fF
C22 VREF m1_688_1652# 0.23fF
C23 INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# VDD 1.57fF
C24 NMOS_S_74334133_X2_Y1_1679758484_0/a_200_252# m1_688_1652# 0.22fF
C25 VIN STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# 0.00fF
C26 m1_688_1652# m1_2720_1484# 0.00fF
C27 VBIAS m1_688_1652# 0.00fF
C28 m1_1172_1316# VIN 0.00fF
C29 VDD m1_602_1568# 4.71fF
C30 m1_2720_1484# OUT 0.06fF
C31 VDD STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# 4.50fF
C32 NMOS_4T_77406006_X2_Y1_1679758483_1/a_200_252# m1_688_1652# 0.22fF
C33 VREF VIN 0.04fF
C34 STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# m1_602_1568# 0.01fF
C35 m1_1172_1316# VDD 4.38fF
C36 m1_1172_1316# m1_602_1568# 1.07fF
C37 VBIAS VIN 0.00fF
C38 INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# m1_2720_1484# 0.71fF
C39 m1_1172_1316# STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# 0.98fF
C40 VIN m1_688_1652# 0.02fF
C41 VIN VSS 0.13fF
C42 VBIAS VSS 0.01fF
C43 OUT VSS 0.08fF
C44 VDD VSS 19.16fF
C45 NMOS_S_74334133_X2_Y1_1679758484_0/a_200_252# VSS 1.47fF
C46 INV_46031338_PG0_0_0_1679758481_0/m1_312_1400# VSS 1.32fF
C47 NMOS_4T_77406006_X2_Y1_1679758483_1/a_200_252# VSS 1.16fF 
C48 m1_688_1652# VSS 2.23fF
C49 VREF VSS 1.18fF
C50 m1_1172_1316# VSS 0.69fF
C51 m1_2720_1484# VSS 2.76fF
C52 STAGE2_INV_90501218_PG0_0_0_1679758482_0/li_663_571# VSS 2.16fF
.ends
x1 VDD VSS VBIAS VIN VREF OUT comparator
V1 VDD VSS 1.8
V2 VREF VSS 1.5
V3 VBIAS VSS 1.3
V4 VIN VSS sine(0 1.8 100000000)

.tran 10p 100n
.control
run
plot v(VREF) v(VIN) v(VBIAS) V(OUT)
.saveall
.endc
