MACRO TWO_BIT_RES_ADC
  ORIGIN 0 0 ;
  FOREIGN TWO_BIT_RES_ADC 0 0 ;
  SIZE 28.51 BY 45.95 ;
  PIN BIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
      LAYER M2 ;
        RECT 9.72 17.92 10.92 18.2 ;
      LAYER M2 ;
        RECT 9.72 42.28 10.92 42.56 ;
      LAYER M2 ;
        RECT 9.73 2.8 10.05 3.08 ;
      LAYER M3 ;
        RECT 9.75 2.94 10.03 18.06 ;
      LAYER M2 ;
        RECT 9.73 17.92 10.05 18.2 ;
      LAYER M3 ;
        RECT 9.75 18.06 10.03 42.42 ;
      LAYER M2 ;
        RECT 9.73 42.28 10.05 42.56 ;
    END
  END BIAS
  PIN INN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 14.02 12.04 15.22 12.32 ;
      LAYER M2 ;
        RECT 14.02 27.16 15.22 27.44 ;
      LAYER M2 ;
        RECT 14.02 33.04 15.22 33.32 ;
      LAYER M2 ;
        RECT 13.76 12.04 14.19 12.32 ;
      LAYER M3 ;
        RECT 13.62 12.18 13.9 27.3 ;
      LAYER M2 ;
        RECT 13.76 27.16 14.19 27.44 ;
      LAYER M2 ;
        RECT 14.46 27.16 14.78 27.44 ;
      LAYER M1 ;
        RECT 14.495 27.3 14.745 33.18 ;
      LAYER M2 ;
        RECT 14.46 33.04 14.78 33.32 ;
    END
  END INN
  PIN C3
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 25.2 7 26.4 7.28 ;
      LAYER M2 ;
        RECT 25.2 7.84 26.4 8.12 ;
      LAYER M2 ;
        RECT 25.64 7 25.96 7.28 ;
      LAYER M3 ;
        RECT 25.66 7.14 25.94 7.98 ;
      LAYER M2 ;
        RECT 25.64 7.84 25.96 8.12 ;
    END
  END C3
  PIN C2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 25.2 22.12 26.4 22.4 ;
      LAYER M2 ;
        RECT 25.2 22.96 26.4 23.24 ;
      LAYER M2 ;
        RECT 25.64 22.12 25.96 22.4 ;
      LAYER M3 ;
        RECT 25.66 22.26 25.94 23.1 ;
      LAYER M2 ;
        RECT 25.64 22.96 25.96 23.24 ;
    END
  END C2
  PIN C1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 25.2 37.24 26.4 37.52 ;
      LAYER M2 ;
        RECT 25.2 38.08 26.4 38.36 ;
      LAYER M2 ;
        RECT 25.64 37.24 25.96 37.52 ;
      LAYER M3 ;
        RECT 25.66 37.38 25.94 38.22 ;
      LAYER M2 ;
        RECT 25.64 38.08 25.96 38.36 ;
    END
  END C1
  PIN INP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 0.695 0.86 8.335 1.66 ;
    END
  END INP
  OBS 
  LAYER M4 ;
        RECT 0.695 9.68 8.335 10.48 ;
  LAYER M4 ;
        RECT 0.695 12.2 8.335 13 ;
  LAYER M4 ;
        RECT 4.275 9.68 4.605 10.48 ;
  LAYER M5 ;
        RECT 3.85 10.08 5.03 12.6 ;
  LAYER M4 ;
        RECT 4.275 12.2 4.605 13 ;
  LAYER M2 ;
        RECT 10.58 12.04 11.78 12.32 ;
  LAYER M4 ;
        RECT 8.005 12.2 8.335 13 ;
  LAYER M3 ;
        RECT 8.03 12.18 8.31 12.6 ;
  LAYER M2 ;
        RECT 8.17 12.04 10.75 12.32 ;
  LAYER M2 ;
        RECT 8.01 12.04 8.33 12.32 ;
  LAYER M3 ;
        RECT 8.03 12.02 8.31 12.34 ;
  LAYER M3 ;
        RECT 8.03 12.415 8.31 12.785 ;
  LAYER M4 ;
        RECT 8.005 12.2 8.335 13 ;
  LAYER M2 ;
        RECT 8.01 12.04 8.33 12.32 ;
  LAYER M3 ;
        RECT 8.03 12.02 8.31 12.34 ;
  LAYER M3 ;
        RECT 8.03 12.415 8.31 12.785 ;
  LAYER M4 ;
        RECT 8.005 12.2 8.335 13 ;
  LAYER M4 ;
        RECT 0.695 21.02 8.335 21.82 ;
  LAYER M4 ;
        RECT 0.695 23.54 8.335 24.34 ;
  LAYER M2 ;
        RECT 10.58 27.16 11.78 27.44 ;
  LAYER M4 ;
        RECT 6.715 21.02 7.045 21.82 ;
  LAYER M3 ;
        RECT 6.74 21.42 7.02 23.94 ;
  LAYER M4 ;
        RECT 6.715 23.54 7.045 24.34 ;
  LAYER M4 ;
        RECT 8.005 23.54 8.335 24.34 ;
  LAYER M3 ;
        RECT 8.03 23.94 8.31 27.3 ;
  LAYER M2 ;
        RECT 8.17 27.16 10.75 27.44 ;
  LAYER M3 ;
        RECT 6.74 21.235 7.02 21.605 ;
  LAYER M4 ;
        RECT 6.715 21.02 7.045 21.82 ;
  LAYER M3 ;
        RECT 6.74 23.755 7.02 24.125 ;
  LAYER M4 ;
        RECT 6.715 23.54 7.045 24.34 ;
  LAYER M3 ;
        RECT 6.74 21.235 7.02 21.605 ;
  LAYER M4 ;
        RECT 6.715 21.02 7.045 21.82 ;
  LAYER M3 ;
        RECT 6.74 23.755 7.02 24.125 ;
  LAYER M4 ;
        RECT 6.715 23.54 7.045 24.34 ;
  LAYER M2 ;
        RECT 8.01 27.16 8.33 27.44 ;
  LAYER M3 ;
        RECT 8.03 27.14 8.31 27.46 ;
  LAYER M3 ;
        RECT 6.74 21.235 7.02 21.605 ;
  LAYER M4 ;
        RECT 6.715 21.02 7.045 21.82 ;
  LAYER M3 ;
        RECT 6.74 23.755 7.02 24.125 ;
  LAYER M4 ;
        RECT 6.715 23.54 7.045 24.34 ;
  LAYER M3 ;
        RECT 8.03 23.755 8.31 24.125 ;
  LAYER M4 ;
        RECT 8.005 23.54 8.335 24.34 ;
  LAYER M2 ;
        RECT 8.01 27.16 8.33 27.44 ;
  LAYER M3 ;
        RECT 8.03 27.14 8.31 27.46 ;
  LAYER M3 ;
        RECT 6.74 21.235 7.02 21.605 ;
  LAYER M4 ;
        RECT 6.715 21.02 7.045 21.82 ;
  LAYER M3 ;
        RECT 6.74 23.755 7.02 24.125 ;
  LAYER M4 ;
        RECT 6.715 23.54 7.045 24.34 ;
  LAYER M3 ;
        RECT 8.03 23.755 8.31 24.125 ;
  LAYER M4 ;
        RECT 8.005 23.54 8.335 24.34 ;
  LAYER M4 ;
        RECT 0.695 32.36 8.335 33.16 ;
  LAYER M4 ;
        RECT 0.695 34.88 8.335 35.68 ;
  LAYER M4 ;
        RECT 4.275 32.36 4.605 33.16 ;
  LAYER M5 ;
        RECT 3.85 32.76 5.03 35.28 ;
  LAYER M4 ;
        RECT 4.275 34.88 4.605 35.68 ;
  LAYER M2 ;
        RECT 10.58 33.04 11.78 33.32 ;
  LAYER M4 ;
        RECT 8.005 32.36 8.335 33.16 ;
  LAYER M3 ;
        RECT 8.03 32.76 8.31 33.18 ;
  LAYER M2 ;
        RECT 8.17 33.04 10.75 33.32 ;
  LAYER M2 ;
        RECT 8.01 33.04 8.33 33.32 ;
  LAYER M3 ;
        RECT 8.03 33.02 8.31 33.34 ;
  LAYER M3 ;
        RECT 8.03 32.575 8.31 32.945 ;
  LAYER M4 ;
        RECT 8.005 32.36 8.335 33.16 ;
  LAYER M2 ;
        RECT 8.01 33.04 8.33 33.32 ;
  LAYER M3 ;
        RECT 8.03 33.02 8.31 33.34 ;
  LAYER M3 ;
        RECT 8.03 32.575 8.31 32.945 ;
  LAYER M4 ;
        RECT 8.005 32.36 8.335 33.16 ;
  LAYER M2 ;
        RECT 14.02 6.58 15.22 6.86 ;
  LAYER M2 ;
        RECT 14.02 7.84 15.22 8.12 ;
  LAYER M2 ;
        RECT 18.32 2.8 19.52 3.08 ;
  LAYER M2 ;
        RECT 18.32 12.04 19.52 12.32 ;
  LAYER M2 ;
        RECT 18.76 2.8 19.08 3.08 ;
  LAYER M3 ;
        RECT 18.78 2.94 19.06 12.18 ;
  LAYER M2 ;
        RECT 18.76 12.04 19.08 12.32 ;
  LAYER M2 ;
        RECT 14.46 6.58 14.78 6.86 ;
  LAYER M3 ;
        RECT 14.48 6.72 14.76 7.98 ;
  LAYER M2 ;
        RECT 14.46 7.84 14.78 8.12 ;
  LAYER M3 ;
        RECT 14.48 7.375 14.76 7.745 ;
  LAYER M2 ;
        RECT 14.62 7.42 18.92 7.7 ;
  LAYER M3 ;
        RECT 18.78 7.375 19.06 7.745 ;
  LAYER M2 ;
        RECT 14.46 6.58 14.78 6.86 ;
  LAYER M3 ;
        RECT 14.48 6.56 14.76 6.88 ;
  LAYER M2 ;
        RECT 14.46 7.84 14.78 8.12 ;
  LAYER M3 ;
        RECT 14.48 7.82 14.76 8.14 ;
  LAYER M2 ;
        RECT 14.46 6.58 14.78 6.86 ;
  LAYER M3 ;
        RECT 14.48 6.56 14.76 6.88 ;
  LAYER M2 ;
        RECT 14.46 7.84 14.78 8.12 ;
  LAYER M3 ;
        RECT 14.48 7.82 14.76 8.14 ;
  LAYER M2 ;
        RECT 14.46 6.58 14.78 6.86 ;
  LAYER M3 ;
        RECT 14.48 6.56 14.76 6.88 ;
  LAYER M2 ;
        RECT 14.46 7.42 14.78 7.7 ;
  LAYER M3 ;
        RECT 14.48 7.4 14.76 7.72 ;
  LAYER M2 ;
        RECT 14.46 7.84 14.78 8.12 ;
  LAYER M3 ;
        RECT 14.48 7.82 14.76 8.14 ;
  LAYER M2 ;
        RECT 18.76 7.42 19.08 7.7 ;
  LAYER M3 ;
        RECT 18.78 7.4 19.06 7.72 ;
  LAYER M2 ;
        RECT 14.46 6.58 14.78 6.86 ;
  LAYER M3 ;
        RECT 14.48 6.56 14.76 6.88 ;
  LAYER M2 ;
        RECT 14.46 7.42 14.78 7.7 ;
  LAYER M3 ;
        RECT 14.48 7.4 14.76 7.72 ;
  LAYER M2 ;
        RECT 14.46 7.84 14.78 8.12 ;
  LAYER M3 ;
        RECT 14.48 7.82 14.76 8.14 ;
  LAYER M2 ;
        RECT 18.76 7.42 19.08 7.7 ;
  LAYER M3 ;
        RECT 18.78 7.4 19.06 7.72 ;
  LAYER M2 ;
        RECT 25.2 2.8 26.4 3.08 ;
  LAYER M2 ;
        RECT 25.2 12.04 26.4 12.32 ;
  LAYER M2 ;
        RECT 25.21 2.8 25.53 3.08 ;
  LAYER M3 ;
        RECT 25.23 2.94 25.51 12.18 ;
  LAYER M2 ;
        RECT 25.21 12.04 25.53 12.32 ;
  LAYER M2 ;
        RECT 21.76 7 22.96 7.28 ;
  LAYER M2 ;
        RECT 21.76 7.84 22.96 8.12 ;
  LAYER M2 ;
        RECT 22.2 7 22.52 7.28 ;
  LAYER M3 ;
        RECT 22.22 7.14 22.5 7.98 ;
  LAYER M2 ;
        RECT 22.2 7.84 22.52 8.12 ;
  LAYER M3 ;
        RECT 25.23 7.375 25.51 7.745 ;
  LAYER M2 ;
        RECT 22.36 7.42 25.37 7.7 ;
  LAYER M3 ;
        RECT 22.22 7.375 22.5 7.745 ;
  LAYER M2 ;
        RECT 22.2 7.42 22.52 7.7 ;
  LAYER M3 ;
        RECT 22.22 7.4 22.5 7.72 ;
  LAYER M2 ;
        RECT 25.21 7.42 25.53 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.4 25.51 7.72 ;
  LAYER M2 ;
        RECT 22.2 7.42 22.52 7.7 ;
  LAYER M3 ;
        RECT 22.22 7.4 22.5 7.72 ;
  LAYER M2 ;
        RECT 25.21 7.42 25.53 7.7 ;
  LAYER M3 ;
        RECT 25.23 7.4 25.51 7.72 ;
  LAYER M2 ;
        RECT 10.58 7.84 11.78 8.12 ;
  LAYER M3 ;
        RECT 14.05 2.78 14.33 7.3 ;
  LAYER M2 ;
        RECT 11.61 7.84 12.9 8.12 ;
  LAYER M3 ;
        RECT 12.76 7.56 13.04 7.98 ;
  LAYER M4 ;
        RECT 12.9 7.16 14.19 7.96 ;
  LAYER M3 ;
        RECT 14.05 7.14 14.33 7.56 ;
  LAYER M2 ;
        RECT 12.74 7.84 13.06 8.12 ;
  LAYER M3 ;
        RECT 12.76 7.82 13.04 8.14 ;
  LAYER M3 ;
        RECT 12.76 7.375 13.04 7.745 ;
  LAYER M4 ;
        RECT 12.735 7.16 13.065 7.96 ;
  LAYER M3 ;
        RECT 14.05 7.375 14.33 7.745 ;
  LAYER M4 ;
        RECT 14.025 7.16 14.355 7.96 ;
  LAYER M2 ;
        RECT 12.74 7.84 13.06 8.12 ;
  LAYER M3 ;
        RECT 12.76 7.82 13.04 8.14 ;
  LAYER M3 ;
        RECT 12.76 7.375 13.04 7.745 ;
  LAYER M4 ;
        RECT 12.735 7.16 13.065 7.96 ;
  LAYER M3 ;
        RECT 14.05 7.375 14.33 7.745 ;
  LAYER M4 ;
        RECT 14.025 7.16 14.355 7.96 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 10.15 8.26 12.21 8.54 ;
  LAYER M2 ;
        RECT 13.59 8.26 15.65 8.54 ;
  LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
  LAYER M3 ;
        RECT 10.18 7.14 10.46 8.4 ;
  LAYER M2 ;
        RECT 10.16 8.26 10.48 8.54 ;
  LAYER M2 ;
        RECT 12.04 8.26 13.76 8.54 ;
  LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
  LAYER M3 ;
        RECT 10.18 6.98 10.46 7.3 ;
  LAYER M2 ;
        RECT 10.16 8.26 10.48 8.54 ;
  LAYER M3 ;
        RECT 10.18 8.24 10.46 8.56 ;
  LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
  LAYER M3 ;
        RECT 10.18 6.98 10.46 7.3 ;
  LAYER M2 ;
        RECT 10.16 8.26 10.48 8.54 ;
  LAYER M3 ;
        RECT 10.18 8.24 10.46 8.56 ;
  LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
  LAYER M3 ;
        RECT 10.18 6.98 10.46 7.3 ;
  LAYER M2 ;
        RECT 10.16 8.26 10.48 8.54 ;
  LAYER M3 ;
        RECT 10.18 8.24 10.46 8.56 ;
  LAYER M2 ;
        RECT 10.16 7 10.48 7.28 ;
  LAYER M3 ;
        RECT 10.18 6.98 10.46 7.3 ;
  LAYER M2 ;
        RECT 10.16 8.26 10.48 8.54 ;
  LAYER M3 ;
        RECT 10.18 8.24 10.46 8.56 ;
  LAYER M2 ;
        RECT 21.76 2.8 22.96 3.08 ;
  LAYER M2 ;
        RECT 18.32 7 19.52 7.28 ;
  LAYER M2 ;
        RECT 18.32 7.84 19.52 8.12 ;
  LAYER M2 ;
        RECT 21.76 12.04 22.96 12.32 ;
  LAYER M2 ;
        RECT 20.64 2.8 21.93 3.08 ;
  LAYER M1 ;
        RECT 20.515 2.94 20.765 7.14 ;
  LAYER M2 ;
        RECT 19.35 7 20.64 7.28 ;
  LAYER M2 ;
        RECT 19.19 7 19.51 7.28 ;
  LAYER M3 ;
        RECT 19.21 7.14 19.49 7.98 ;
  LAYER M2 ;
        RECT 19.19 7.84 19.51 8.12 ;
  LAYER M1 ;
        RECT 20.515 7.14 20.765 12.18 ;
  LAYER M2 ;
        RECT 20.64 12.04 21.93 12.32 ;
  LAYER M1 ;
        RECT 20.515 2.855 20.765 3.025 ;
  LAYER M2 ;
        RECT 20.47 2.8 20.81 3.08 ;
  LAYER M1 ;
        RECT 20.515 7.055 20.765 7.225 ;
  LAYER M2 ;
        RECT 20.47 7 20.81 7.28 ;
  LAYER M1 ;
        RECT 20.515 2.855 20.765 3.025 ;
  LAYER M2 ;
        RECT 20.47 2.8 20.81 3.08 ;
  LAYER M1 ;
        RECT 20.515 7.055 20.765 7.225 ;
  LAYER M2 ;
        RECT 20.47 7 20.81 7.28 ;
  LAYER M1 ;
        RECT 20.515 2.855 20.765 3.025 ;
  LAYER M2 ;
        RECT 20.47 2.8 20.81 3.08 ;
  LAYER M1 ;
        RECT 20.515 7.055 20.765 7.225 ;
  LAYER M2 ;
        RECT 20.47 7 20.81 7.28 ;
  LAYER M2 ;
        RECT 19.19 7 19.51 7.28 ;
  LAYER M3 ;
        RECT 19.21 6.98 19.49 7.3 ;
  LAYER M2 ;
        RECT 19.19 7.84 19.51 8.12 ;
  LAYER M3 ;
        RECT 19.21 7.82 19.49 8.14 ;
  LAYER M1 ;
        RECT 20.515 2.855 20.765 3.025 ;
  LAYER M2 ;
        RECT 20.47 2.8 20.81 3.08 ;
  LAYER M1 ;
        RECT 20.515 7.055 20.765 7.225 ;
  LAYER M2 ;
        RECT 20.47 7 20.81 7.28 ;
  LAYER M2 ;
        RECT 19.19 7 19.51 7.28 ;
  LAYER M3 ;
        RECT 19.21 6.98 19.49 7.3 ;
  LAYER M2 ;
        RECT 19.19 7.84 19.51 8.12 ;
  LAYER M3 ;
        RECT 19.21 7.82 19.49 8.14 ;
  LAYER M1 ;
        RECT 20.515 2.855 20.765 3.025 ;
  LAYER M2 ;
        RECT 20.47 2.8 20.81 3.08 ;
  LAYER M1 ;
        RECT 20.515 7.055 20.765 7.225 ;
  LAYER M2 ;
        RECT 20.47 7 20.81 7.28 ;
  LAYER M1 ;
        RECT 20.515 12.095 20.765 12.265 ;
  LAYER M2 ;
        RECT 20.47 12.04 20.81 12.32 ;
  LAYER M2 ;
        RECT 19.19 7 19.51 7.28 ;
  LAYER M3 ;
        RECT 19.21 6.98 19.49 7.3 ;
  LAYER M2 ;
        RECT 19.19 7.84 19.51 8.12 ;
  LAYER M3 ;
        RECT 19.21 7.82 19.49 8.14 ;
  LAYER M1 ;
        RECT 20.515 2.855 20.765 3.025 ;
  LAYER M2 ;
        RECT 20.47 2.8 20.81 3.08 ;
  LAYER M1 ;
        RECT 20.515 7.055 20.765 7.225 ;
  LAYER M2 ;
        RECT 20.47 7 20.81 7.28 ;
  LAYER M1 ;
        RECT 20.515 12.095 20.765 12.265 ;
  LAYER M2 ;
        RECT 20.47 12.04 20.81 12.32 ;
  LAYER M2 ;
        RECT 19.19 7 19.51 7.28 ;
  LAYER M3 ;
        RECT 19.21 6.98 19.49 7.3 ;
  LAYER M2 ;
        RECT 19.19 7.84 19.51 8.12 ;
  LAYER M3 ;
        RECT 19.21 7.82 19.49 8.14 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 18.365 3.695 18.615 7.225 ;
  LAYER M1 ;
        RECT 18.365 2.435 18.615 3.445 ;
  LAYER M1 ;
        RECT 18.365 0.335 18.615 1.345 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M2 ;
        RECT 17.89 6.58 19.95 6.86 ;
  LAYER M2 ;
        RECT 18.32 0.7 19.52 0.98 ;
  LAYER M2 ;
        RECT 18.32 7 19.52 7.28 ;
  LAYER M2 ;
        RECT 18.32 2.8 19.52 3.08 ;
  LAYER M3 ;
        RECT 18.35 0.68 18.63 6.88 ;
  LAYER M1 ;
        RECT 22.665 3.695 22.915 7.225 ;
  LAYER M1 ;
        RECT 22.665 2.435 22.915 3.445 ;
  LAYER M1 ;
        RECT 22.665 0.335 22.915 1.345 ;
  LAYER M1 ;
        RECT 23.095 3.695 23.345 7.225 ;
  LAYER M1 ;
        RECT 22.235 3.695 22.485 7.225 ;
  LAYER M1 ;
        RECT 21.805 3.695 22.055 7.225 ;
  LAYER M1 ;
        RECT 21.805 2.435 22.055 3.445 ;
  LAYER M1 ;
        RECT 21.805 0.335 22.055 1.345 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M2 ;
        RECT 21.33 6.58 23.39 6.86 ;
  LAYER M2 ;
        RECT 21.76 0.7 22.96 0.98 ;
  LAYER M2 ;
        RECT 21.76 7 22.96 7.28 ;
  LAYER M2 ;
        RECT 21.76 2.8 22.96 3.08 ;
  LAYER M3 ;
        RECT 21.79 0.68 22.07 6.88 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 11.425 ;
  LAYER M1 ;
        RECT 19.225 11.675 19.475 12.685 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 14.785 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M1 ;
        RECT 18.795 7.895 19.045 11.425 ;
  LAYER M1 ;
        RECT 18.365 7.895 18.615 11.425 ;
  LAYER M1 ;
        RECT 18.365 11.675 18.615 12.685 ;
  LAYER M1 ;
        RECT 18.365 13.775 18.615 14.785 ;
  LAYER M1 ;
        RECT 17.935 7.895 18.185 11.425 ;
  LAYER M2 ;
        RECT 17.89 8.26 19.95 8.54 ;
  LAYER M2 ;
        RECT 18.32 14.14 19.52 14.42 ;
  LAYER M2 ;
        RECT 18.32 7.84 19.52 8.12 ;
  LAYER M2 ;
        RECT 18.32 12.04 19.52 12.32 ;
  LAYER M3 ;
        RECT 18.35 8.24 18.63 14.44 ;
  LAYER M1 ;
        RECT 22.665 7.895 22.915 11.425 ;
  LAYER M1 ;
        RECT 22.665 11.675 22.915 12.685 ;
  LAYER M1 ;
        RECT 22.665 13.775 22.915 14.785 ;
  LAYER M1 ;
        RECT 23.095 7.895 23.345 11.425 ;
  LAYER M1 ;
        RECT 22.235 7.895 22.485 11.425 ;
  LAYER M1 ;
        RECT 21.805 7.895 22.055 11.425 ;
  LAYER M1 ;
        RECT 21.805 11.675 22.055 12.685 ;
  LAYER M1 ;
        RECT 21.805 13.775 22.055 14.785 ;
  LAYER M1 ;
        RECT 21.375 7.895 21.625 11.425 ;
  LAYER M2 ;
        RECT 21.33 8.26 23.39 8.54 ;
  LAYER M2 ;
        RECT 21.76 14.14 22.96 14.42 ;
  LAYER M2 ;
        RECT 21.76 7.84 22.96 8.12 ;
  LAYER M2 ;
        RECT 21.76 12.04 22.96 12.32 ;
  LAYER M3 ;
        RECT 21.79 8.24 22.07 14.44 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M1 ;
        RECT 15.785 3.695 16.035 7.225 ;
  LAYER M1 ;
        RECT 15.785 2.435 16.035 3.445 ;
  LAYER M1 ;
        RECT 15.785 0.335 16.035 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M2 ;
        RECT 13.16 7 16.08 7.28 ;
  LAYER M2 ;
        RECT 13.16 2.8 16.08 3.08 ;
  LAYER M2 ;
        RECT 12.73 6.16 16.51 6.44 ;
  LAYER M2 ;
        RECT 13.16 0.7 16.08 0.98 ;
  LAYER M3 ;
        RECT 14.05 2.78 14.33 7.3 ;
  LAYER M2 ;
        RECT 14.02 6.58 15.22 6.86 ;
  LAYER M3 ;
        RECT 14.91 0.68 15.19 6.46 ;
  LAYER M1 ;
        RECT 25.245 3.695 25.495 7.225 ;
  LAYER M1 ;
        RECT 25.245 2.435 25.495 3.445 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 1.345 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M1 ;
        RECT 25.675 3.695 25.925 7.225 ;
  LAYER M1 ;
        RECT 26.105 3.695 26.355 7.225 ;
  LAYER M1 ;
        RECT 26.105 2.435 26.355 3.445 ;
  LAYER M1 ;
        RECT 26.105 0.335 26.355 1.345 ;
  LAYER M1 ;
        RECT 26.535 3.695 26.785 7.225 ;
  LAYER M2 ;
        RECT 24.77 6.58 26.83 6.86 ;
  LAYER M2 ;
        RECT 25.2 0.7 26.4 0.98 ;
  LAYER M2 ;
        RECT 25.2 7 26.4 7.28 ;
  LAYER M2 ;
        RECT 25.2 2.8 26.4 3.08 ;
  LAYER M3 ;
        RECT 26.09 0.68 26.37 6.88 ;
  LAYER M1 ;
        RECT 25.245 7.895 25.495 11.425 ;
  LAYER M1 ;
        RECT 25.245 11.675 25.495 12.685 ;
  LAYER M1 ;
        RECT 25.245 13.775 25.495 14.785 ;
  LAYER M1 ;
        RECT 24.815 7.895 25.065 11.425 ;
  LAYER M1 ;
        RECT 25.675 7.895 25.925 11.425 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 11.425 ;
  LAYER M1 ;
        RECT 26.105 11.675 26.355 12.685 ;
  LAYER M1 ;
        RECT 26.105 13.775 26.355 14.785 ;
  LAYER M1 ;
        RECT 26.535 7.895 26.785 11.425 ;
  LAYER M2 ;
        RECT 24.77 8.26 26.83 8.54 ;
  LAYER M2 ;
        RECT 25.2 14.14 26.4 14.42 ;
  LAYER M2 ;
        RECT 25.2 7.84 26.4 8.12 ;
  LAYER M2 ;
        RECT 25.2 12.04 26.4 12.32 ;
  LAYER M3 ;
        RECT 26.09 8.24 26.37 14.44 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M2 ;
        RECT 9.29 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 9.72 0.7 10.92 0.98 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M3 ;
        RECT 10.61 0.68 10.89 6.88 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M2 ;
        RECT 10.58 14.14 11.78 14.42 ;
  LAYER M2 ;
        RECT 10.58 7.84 11.78 8.12 ;
  LAYER M2 ;
        RECT 10.58 12.04 11.78 12.32 ;
  LAYER M2 ;
        RECT 10.15 8.26 12.21 8.54 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 11.425 ;
  LAYER M1 ;
        RECT 14.925 11.675 15.175 12.685 ;
  LAYER M1 ;
        RECT 14.925 13.775 15.175 14.785 ;
  LAYER M1 ;
        RECT 15.355 7.895 15.605 11.425 ;
  LAYER M2 ;
        RECT 14.02 14.14 15.22 14.42 ;
  LAYER M2 ;
        RECT 14.02 7.84 15.22 8.12 ;
  LAYER M2 ;
        RECT 14.02 12.04 15.22 12.32 ;
  LAYER M2 ;
        RECT 13.59 8.26 15.65 8.54 ;
  LAYER M2 ;
        RECT 14.02 21.7 15.22 21.98 ;
  LAYER M2 ;
        RECT 14.02 22.96 15.22 23.24 ;
  LAYER M2 ;
        RECT 18.32 17.92 19.52 18.2 ;
  LAYER M2 ;
        RECT 18.32 27.16 19.52 27.44 ;
  LAYER M2 ;
        RECT 18.76 17.92 19.08 18.2 ;
  LAYER M3 ;
        RECT 18.78 18.06 19.06 27.3 ;
  LAYER M2 ;
        RECT 18.76 27.16 19.08 27.44 ;
  LAYER M2 ;
        RECT 14.46 21.7 14.78 21.98 ;
  LAYER M3 ;
        RECT 14.48 21.84 14.76 23.1 ;
  LAYER M2 ;
        RECT 14.46 22.96 14.78 23.24 ;
  LAYER M3 ;
        RECT 14.48 22.495 14.76 22.865 ;
  LAYER M2 ;
        RECT 14.62 22.54 18.92 22.82 ;
  LAYER M3 ;
        RECT 18.78 22.495 19.06 22.865 ;
  LAYER M2 ;
        RECT 14.46 21.7 14.78 21.98 ;
  LAYER M3 ;
        RECT 14.48 21.68 14.76 22 ;
  LAYER M2 ;
        RECT 14.46 22.96 14.78 23.24 ;
  LAYER M3 ;
        RECT 14.48 22.94 14.76 23.26 ;
  LAYER M2 ;
        RECT 14.46 21.7 14.78 21.98 ;
  LAYER M3 ;
        RECT 14.48 21.68 14.76 22 ;
  LAYER M2 ;
        RECT 14.46 22.96 14.78 23.24 ;
  LAYER M3 ;
        RECT 14.48 22.94 14.76 23.26 ;
  LAYER M2 ;
        RECT 14.46 21.7 14.78 21.98 ;
  LAYER M3 ;
        RECT 14.48 21.68 14.76 22 ;
  LAYER M2 ;
        RECT 14.46 22.54 14.78 22.82 ;
  LAYER M3 ;
        RECT 14.48 22.52 14.76 22.84 ;
  LAYER M2 ;
        RECT 14.46 22.96 14.78 23.24 ;
  LAYER M3 ;
        RECT 14.48 22.94 14.76 23.26 ;
  LAYER M2 ;
        RECT 18.76 22.54 19.08 22.82 ;
  LAYER M3 ;
        RECT 18.78 22.52 19.06 22.84 ;
  LAYER M2 ;
        RECT 14.46 21.7 14.78 21.98 ;
  LAYER M3 ;
        RECT 14.48 21.68 14.76 22 ;
  LAYER M2 ;
        RECT 14.46 22.54 14.78 22.82 ;
  LAYER M3 ;
        RECT 14.48 22.52 14.76 22.84 ;
  LAYER M2 ;
        RECT 14.46 22.96 14.78 23.24 ;
  LAYER M3 ;
        RECT 14.48 22.94 14.76 23.26 ;
  LAYER M2 ;
        RECT 18.76 22.54 19.08 22.82 ;
  LAYER M3 ;
        RECT 18.78 22.52 19.06 22.84 ;
  LAYER M2 ;
        RECT 25.2 17.92 26.4 18.2 ;
  LAYER M2 ;
        RECT 25.2 27.16 26.4 27.44 ;
  LAYER M2 ;
        RECT 25.21 17.92 25.53 18.2 ;
  LAYER M3 ;
        RECT 25.23 18.06 25.51 27.3 ;
  LAYER M2 ;
        RECT 25.21 27.16 25.53 27.44 ;
  LAYER M2 ;
        RECT 21.76 22.12 22.96 22.4 ;
  LAYER M2 ;
        RECT 21.76 22.96 22.96 23.24 ;
  LAYER M2 ;
        RECT 22.2 22.12 22.52 22.4 ;
  LAYER M3 ;
        RECT 22.22 22.26 22.5 23.1 ;
  LAYER M2 ;
        RECT 22.2 22.96 22.52 23.24 ;
  LAYER M3 ;
        RECT 25.23 22.495 25.51 22.865 ;
  LAYER M2 ;
        RECT 22.36 22.54 25.37 22.82 ;
  LAYER M3 ;
        RECT 22.22 22.495 22.5 22.865 ;
  LAYER M2 ;
        RECT 22.2 22.54 22.52 22.82 ;
  LAYER M3 ;
        RECT 22.22 22.52 22.5 22.84 ;
  LAYER M2 ;
        RECT 25.21 22.54 25.53 22.82 ;
  LAYER M3 ;
        RECT 25.23 22.52 25.51 22.84 ;
  LAYER M2 ;
        RECT 22.2 22.54 22.52 22.82 ;
  LAYER M3 ;
        RECT 22.22 22.52 22.5 22.84 ;
  LAYER M2 ;
        RECT 25.21 22.54 25.53 22.82 ;
  LAYER M3 ;
        RECT 25.23 22.52 25.51 22.84 ;
  LAYER M2 ;
        RECT 10.58 22.96 11.78 23.24 ;
  LAYER M3 ;
        RECT 14.05 17.9 14.33 22.42 ;
  LAYER M2 ;
        RECT 11.61 22.96 13.33 23.24 ;
  LAYER M3 ;
        RECT 13.19 22.68 13.47 23.1 ;
  LAYER M4 ;
        RECT 13.33 22.28 14.19 23.08 ;
  LAYER M3 ;
        RECT 14.05 22.26 14.33 22.68 ;
  LAYER M2 ;
        RECT 13.17 22.96 13.49 23.24 ;
  LAYER M3 ;
        RECT 13.19 22.94 13.47 23.26 ;
  LAYER M3 ;
        RECT 13.19 22.495 13.47 22.865 ;
  LAYER M4 ;
        RECT 13.165 22.28 13.495 23.08 ;
  LAYER M3 ;
        RECT 14.05 22.495 14.33 22.865 ;
  LAYER M4 ;
        RECT 14.025 22.28 14.355 23.08 ;
  LAYER M2 ;
        RECT 13.17 22.96 13.49 23.24 ;
  LAYER M3 ;
        RECT 13.19 22.94 13.47 23.26 ;
  LAYER M3 ;
        RECT 13.19 22.495 13.47 22.865 ;
  LAYER M4 ;
        RECT 13.165 22.28 13.495 23.08 ;
  LAYER M3 ;
        RECT 14.05 22.495 14.33 22.865 ;
  LAYER M4 ;
        RECT 14.025 22.28 14.355 23.08 ;
  LAYER M2 ;
        RECT 9.72 22.12 10.92 22.4 ;
  LAYER M2 ;
        RECT 10.15 23.38 12.21 23.66 ;
  LAYER M2 ;
        RECT 13.59 23.38 15.65 23.66 ;
  LAYER M2 ;
        RECT 10.16 22.12 10.48 22.4 ;
  LAYER M3 ;
        RECT 10.18 22.26 10.46 23.52 ;
  LAYER M2 ;
        RECT 10.16 23.38 10.48 23.66 ;
  LAYER M2 ;
        RECT 12.04 23.38 13.76 23.66 ;
  LAYER M2 ;
        RECT 10.16 22.12 10.48 22.4 ;
  LAYER M3 ;
        RECT 10.18 22.1 10.46 22.42 ;
  LAYER M2 ;
        RECT 10.16 23.38 10.48 23.66 ;
  LAYER M3 ;
        RECT 10.18 23.36 10.46 23.68 ;
  LAYER M2 ;
        RECT 10.16 22.12 10.48 22.4 ;
  LAYER M3 ;
        RECT 10.18 22.1 10.46 22.42 ;
  LAYER M2 ;
        RECT 10.16 23.38 10.48 23.66 ;
  LAYER M3 ;
        RECT 10.18 23.36 10.46 23.68 ;
  LAYER M2 ;
        RECT 10.16 22.12 10.48 22.4 ;
  LAYER M3 ;
        RECT 10.18 22.1 10.46 22.42 ;
  LAYER M2 ;
        RECT 10.16 23.38 10.48 23.66 ;
  LAYER M3 ;
        RECT 10.18 23.36 10.46 23.68 ;
  LAYER M2 ;
        RECT 10.16 22.12 10.48 22.4 ;
  LAYER M3 ;
        RECT 10.18 22.1 10.46 22.42 ;
  LAYER M2 ;
        RECT 10.16 23.38 10.48 23.66 ;
  LAYER M3 ;
        RECT 10.18 23.36 10.46 23.68 ;
  LAYER M2 ;
        RECT 21.76 17.92 22.96 18.2 ;
  LAYER M2 ;
        RECT 18.32 22.12 19.52 22.4 ;
  LAYER M2 ;
        RECT 18.32 22.96 19.52 23.24 ;
  LAYER M2 ;
        RECT 21.76 27.16 22.96 27.44 ;
  LAYER M2 ;
        RECT 20.64 17.92 21.93 18.2 ;
  LAYER M1 ;
        RECT 20.515 18.06 20.765 22.26 ;
  LAYER M2 ;
        RECT 19.35 22.12 20.64 22.4 ;
  LAYER M2 ;
        RECT 19.19 22.12 19.51 22.4 ;
  LAYER M3 ;
        RECT 19.21 22.26 19.49 23.1 ;
  LAYER M2 ;
        RECT 19.19 22.96 19.51 23.24 ;
  LAYER M1 ;
        RECT 20.515 22.26 20.765 27.3 ;
  LAYER M2 ;
        RECT 20.64 27.16 21.93 27.44 ;
  LAYER M1 ;
        RECT 20.515 17.975 20.765 18.145 ;
  LAYER M2 ;
        RECT 20.47 17.92 20.81 18.2 ;
  LAYER M1 ;
        RECT 20.515 22.175 20.765 22.345 ;
  LAYER M2 ;
        RECT 20.47 22.12 20.81 22.4 ;
  LAYER M1 ;
        RECT 20.515 17.975 20.765 18.145 ;
  LAYER M2 ;
        RECT 20.47 17.92 20.81 18.2 ;
  LAYER M1 ;
        RECT 20.515 22.175 20.765 22.345 ;
  LAYER M2 ;
        RECT 20.47 22.12 20.81 22.4 ;
  LAYER M1 ;
        RECT 20.515 17.975 20.765 18.145 ;
  LAYER M2 ;
        RECT 20.47 17.92 20.81 18.2 ;
  LAYER M1 ;
        RECT 20.515 22.175 20.765 22.345 ;
  LAYER M2 ;
        RECT 20.47 22.12 20.81 22.4 ;
  LAYER M2 ;
        RECT 19.19 22.12 19.51 22.4 ;
  LAYER M3 ;
        RECT 19.21 22.1 19.49 22.42 ;
  LAYER M2 ;
        RECT 19.19 22.96 19.51 23.24 ;
  LAYER M3 ;
        RECT 19.21 22.94 19.49 23.26 ;
  LAYER M1 ;
        RECT 20.515 17.975 20.765 18.145 ;
  LAYER M2 ;
        RECT 20.47 17.92 20.81 18.2 ;
  LAYER M1 ;
        RECT 20.515 22.175 20.765 22.345 ;
  LAYER M2 ;
        RECT 20.47 22.12 20.81 22.4 ;
  LAYER M2 ;
        RECT 19.19 22.12 19.51 22.4 ;
  LAYER M3 ;
        RECT 19.21 22.1 19.49 22.42 ;
  LAYER M2 ;
        RECT 19.19 22.96 19.51 23.24 ;
  LAYER M3 ;
        RECT 19.21 22.94 19.49 23.26 ;
  LAYER M1 ;
        RECT 20.515 17.975 20.765 18.145 ;
  LAYER M2 ;
        RECT 20.47 17.92 20.81 18.2 ;
  LAYER M1 ;
        RECT 20.515 22.175 20.765 22.345 ;
  LAYER M2 ;
        RECT 20.47 22.12 20.81 22.4 ;
  LAYER M1 ;
        RECT 20.515 27.215 20.765 27.385 ;
  LAYER M2 ;
        RECT 20.47 27.16 20.81 27.44 ;
  LAYER M2 ;
        RECT 19.19 22.12 19.51 22.4 ;
  LAYER M3 ;
        RECT 19.21 22.1 19.49 22.42 ;
  LAYER M2 ;
        RECT 19.19 22.96 19.51 23.24 ;
  LAYER M3 ;
        RECT 19.21 22.94 19.49 23.26 ;
  LAYER M1 ;
        RECT 20.515 17.975 20.765 18.145 ;
  LAYER M2 ;
        RECT 20.47 17.92 20.81 18.2 ;
  LAYER M1 ;
        RECT 20.515 22.175 20.765 22.345 ;
  LAYER M2 ;
        RECT 20.47 22.12 20.81 22.4 ;
  LAYER M1 ;
        RECT 20.515 27.215 20.765 27.385 ;
  LAYER M2 ;
        RECT 20.47 27.16 20.81 27.44 ;
  LAYER M2 ;
        RECT 19.19 22.12 19.51 22.4 ;
  LAYER M3 ;
        RECT 19.21 22.1 19.49 22.42 ;
  LAYER M2 ;
        RECT 19.19 22.96 19.51 23.24 ;
  LAYER M3 ;
        RECT 19.21 22.94 19.49 23.26 ;
  LAYER M1 ;
        RECT 19.225 18.815 19.475 22.345 ;
  LAYER M1 ;
        RECT 19.225 17.555 19.475 18.565 ;
  LAYER M1 ;
        RECT 19.225 15.455 19.475 16.465 ;
  LAYER M1 ;
        RECT 19.655 18.815 19.905 22.345 ;
  LAYER M1 ;
        RECT 18.795 18.815 19.045 22.345 ;
  LAYER M1 ;
        RECT 18.365 18.815 18.615 22.345 ;
  LAYER M1 ;
        RECT 18.365 17.555 18.615 18.565 ;
  LAYER M1 ;
        RECT 18.365 15.455 18.615 16.465 ;
  LAYER M1 ;
        RECT 17.935 18.815 18.185 22.345 ;
  LAYER M2 ;
        RECT 17.89 21.7 19.95 21.98 ;
  LAYER M2 ;
        RECT 18.32 15.82 19.52 16.1 ;
  LAYER M2 ;
        RECT 18.32 22.12 19.52 22.4 ;
  LAYER M2 ;
        RECT 18.32 17.92 19.52 18.2 ;
  LAYER M3 ;
        RECT 18.35 15.8 18.63 22 ;
  LAYER M1 ;
        RECT 22.665 18.815 22.915 22.345 ;
  LAYER M1 ;
        RECT 22.665 17.555 22.915 18.565 ;
  LAYER M1 ;
        RECT 22.665 15.455 22.915 16.465 ;
  LAYER M1 ;
        RECT 23.095 18.815 23.345 22.345 ;
  LAYER M1 ;
        RECT 22.235 18.815 22.485 22.345 ;
  LAYER M1 ;
        RECT 21.805 18.815 22.055 22.345 ;
  LAYER M1 ;
        RECT 21.805 17.555 22.055 18.565 ;
  LAYER M1 ;
        RECT 21.805 15.455 22.055 16.465 ;
  LAYER M1 ;
        RECT 21.375 18.815 21.625 22.345 ;
  LAYER M2 ;
        RECT 21.33 21.7 23.39 21.98 ;
  LAYER M2 ;
        RECT 21.76 15.82 22.96 16.1 ;
  LAYER M2 ;
        RECT 21.76 22.12 22.96 22.4 ;
  LAYER M2 ;
        RECT 21.76 17.92 22.96 18.2 ;
  LAYER M3 ;
        RECT 21.79 15.8 22.07 22 ;
  LAYER M1 ;
        RECT 19.225 23.015 19.475 26.545 ;
  LAYER M1 ;
        RECT 19.225 26.795 19.475 27.805 ;
  LAYER M1 ;
        RECT 19.225 28.895 19.475 29.905 ;
  LAYER M1 ;
        RECT 19.655 23.015 19.905 26.545 ;
  LAYER M1 ;
        RECT 18.795 23.015 19.045 26.545 ;
  LAYER M1 ;
        RECT 18.365 23.015 18.615 26.545 ;
  LAYER M1 ;
        RECT 18.365 26.795 18.615 27.805 ;
  LAYER M1 ;
        RECT 18.365 28.895 18.615 29.905 ;
  LAYER M1 ;
        RECT 17.935 23.015 18.185 26.545 ;
  LAYER M2 ;
        RECT 17.89 23.38 19.95 23.66 ;
  LAYER M2 ;
        RECT 18.32 29.26 19.52 29.54 ;
  LAYER M2 ;
        RECT 18.32 22.96 19.52 23.24 ;
  LAYER M2 ;
        RECT 18.32 27.16 19.52 27.44 ;
  LAYER M3 ;
        RECT 18.35 23.36 18.63 29.56 ;
  LAYER M1 ;
        RECT 22.665 23.015 22.915 26.545 ;
  LAYER M1 ;
        RECT 22.665 26.795 22.915 27.805 ;
  LAYER M1 ;
        RECT 22.665 28.895 22.915 29.905 ;
  LAYER M1 ;
        RECT 23.095 23.015 23.345 26.545 ;
  LAYER M1 ;
        RECT 22.235 23.015 22.485 26.545 ;
  LAYER M1 ;
        RECT 21.805 23.015 22.055 26.545 ;
  LAYER M1 ;
        RECT 21.805 26.795 22.055 27.805 ;
  LAYER M1 ;
        RECT 21.805 28.895 22.055 29.905 ;
  LAYER M1 ;
        RECT 21.375 23.015 21.625 26.545 ;
  LAYER M2 ;
        RECT 21.33 23.38 23.39 23.66 ;
  LAYER M2 ;
        RECT 21.76 29.26 22.96 29.54 ;
  LAYER M2 ;
        RECT 21.76 22.96 22.96 23.24 ;
  LAYER M2 ;
        RECT 21.76 27.16 22.96 27.44 ;
  LAYER M3 ;
        RECT 21.79 23.36 22.07 29.56 ;
  LAYER M1 ;
        RECT 13.205 18.815 13.455 22.345 ;
  LAYER M1 ;
        RECT 13.205 17.555 13.455 18.565 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 16.465 ;
  LAYER M1 ;
        RECT 12.775 18.815 13.025 22.345 ;
  LAYER M1 ;
        RECT 13.635 18.815 13.885 22.345 ;
  LAYER M1 ;
        RECT 14.065 18.815 14.315 22.345 ;
  LAYER M1 ;
        RECT 14.065 17.555 14.315 18.565 ;
  LAYER M1 ;
        RECT 14.065 15.455 14.315 16.465 ;
  LAYER M1 ;
        RECT 14.495 18.815 14.745 22.345 ;
  LAYER M1 ;
        RECT 14.925 18.815 15.175 22.345 ;
  LAYER M1 ;
        RECT 14.925 17.555 15.175 18.565 ;
  LAYER M1 ;
        RECT 14.925 15.455 15.175 16.465 ;
  LAYER M1 ;
        RECT 15.355 18.815 15.605 22.345 ;
  LAYER M1 ;
        RECT 15.785 18.815 16.035 22.345 ;
  LAYER M1 ;
        RECT 15.785 17.555 16.035 18.565 ;
  LAYER M1 ;
        RECT 15.785 15.455 16.035 16.465 ;
  LAYER M1 ;
        RECT 16.215 18.815 16.465 22.345 ;
  LAYER M2 ;
        RECT 13.16 22.12 16.08 22.4 ;
  LAYER M2 ;
        RECT 13.16 17.92 16.08 18.2 ;
  LAYER M2 ;
        RECT 12.73 21.28 16.51 21.56 ;
  LAYER M2 ;
        RECT 13.16 15.82 16.08 16.1 ;
  LAYER M3 ;
        RECT 14.05 17.9 14.33 22.42 ;
  LAYER M2 ;
        RECT 14.02 21.7 15.22 21.98 ;
  LAYER M3 ;
        RECT 14.91 15.8 15.19 21.58 ;
  LAYER M1 ;
        RECT 25.245 18.815 25.495 22.345 ;
  LAYER M1 ;
        RECT 25.245 17.555 25.495 18.565 ;
  LAYER M1 ;
        RECT 25.245 15.455 25.495 16.465 ;
  LAYER M1 ;
        RECT 24.815 18.815 25.065 22.345 ;
  LAYER M1 ;
        RECT 25.675 18.815 25.925 22.345 ;
  LAYER M1 ;
        RECT 26.105 18.815 26.355 22.345 ;
  LAYER M1 ;
        RECT 26.105 17.555 26.355 18.565 ;
  LAYER M1 ;
        RECT 26.105 15.455 26.355 16.465 ;
  LAYER M1 ;
        RECT 26.535 18.815 26.785 22.345 ;
  LAYER M2 ;
        RECT 24.77 21.7 26.83 21.98 ;
  LAYER M2 ;
        RECT 25.2 15.82 26.4 16.1 ;
  LAYER M2 ;
        RECT 25.2 22.12 26.4 22.4 ;
  LAYER M2 ;
        RECT 25.2 17.92 26.4 18.2 ;
  LAYER M3 ;
        RECT 26.09 15.8 26.37 22 ;
  LAYER M1 ;
        RECT 25.245 23.015 25.495 26.545 ;
  LAYER M1 ;
        RECT 25.245 26.795 25.495 27.805 ;
  LAYER M1 ;
        RECT 25.245 28.895 25.495 29.905 ;
  LAYER M1 ;
        RECT 24.815 23.015 25.065 26.545 ;
  LAYER M1 ;
        RECT 25.675 23.015 25.925 26.545 ;
  LAYER M1 ;
        RECT 26.105 23.015 26.355 26.545 ;
  LAYER M1 ;
        RECT 26.105 26.795 26.355 27.805 ;
  LAYER M1 ;
        RECT 26.105 28.895 26.355 29.905 ;
  LAYER M1 ;
        RECT 26.535 23.015 26.785 26.545 ;
  LAYER M2 ;
        RECT 24.77 23.38 26.83 23.66 ;
  LAYER M2 ;
        RECT 25.2 29.26 26.4 29.54 ;
  LAYER M2 ;
        RECT 25.2 22.96 26.4 23.24 ;
  LAYER M2 ;
        RECT 25.2 27.16 26.4 27.44 ;
  LAYER M3 ;
        RECT 26.09 23.36 26.37 29.56 ;
  LAYER M1 ;
        RECT 9.765 18.815 10.015 22.345 ;
  LAYER M1 ;
        RECT 9.765 17.555 10.015 18.565 ;
  LAYER M1 ;
        RECT 9.765 15.455 10.015 16.465 ;
  LAYER M1 ;
        RECT 9.335 18.815 9.585 22.345 ;
  LAYER M1 ;
        RECT 10.195 18.815 10.445 22.345 ;
  LAYER M1 ;
        RECT 10.625 18.815 10.875 22.345 ;
  LAYER M1 ;
        RECT 10.625 17.555 10.875 18.565 ;
  LAYER M1 ;
        RECT 10.625 15.455 10.875 16.465 ;
  LAYER M1 ;
        RECT 11.055 18.815 11.305 22.345 ;
  LAYER M2 ;
        RECT 9.29 21.7 11.35 21.98 ;
  LAYER M2 ;
        RECT 9.72 15.82 10.92 16.1 ;
  LAYER M2 ;
        RECT 9.72 22.12 10.92 22.4 ;
  LAYER M2 ;
        RECT 9.72 17.92 10.92 18.2 ;
  LAYER M3 ;
        RECT 10.61 15.8 10.89 22 ;
  LAYER M1 ;
        RECT 10.625 23.015 10.875 26.545 ;
  LAYER M1 ;
        RECT 10.625 26.795 10.875 27.805 ;
  LAYER M1 ;
        RECT 10.625 28.895 10.875 29.905 ;
  LAYER M1 ;
        RECT 10.195 23.015 10.445 26.545 ;
  LAYER M1 ;
        RECT 11.055 23.015 11.305 26.545 ;
  LAYER M1 ;
        RECT 11.485 23.015 11.735 26.545 ;
  LAYER M1 ;
        RECT 11.485 26.795 11.735 27.805 ;
  LAYER M1 ;
        RECT 11.485 28.895 11.735 29.905 ;
  LAYER M1 ;
        RECT 11.915 23.015 12.165 26.545 ;
  LAYER M2 ;
        RECT 10.58 29.26 11.78 29.54 ;
  LAYER M2 ;
        RECT 10.58 22.96 11.78 23.24 ;
  LAYER M2 ;
        RECT 10.58 27.16 11.78 27.44 ;
  LAYER M2 ;
        RECT 10.15 23.38 12.21 23.66 ;
  LAYER M1 ;
        RECT 14.065 23.015 14.315 26.545 ;
  LAYER M1 ;
        RECT 14.065 26.795 14.315 27.805 ;
  LAYER M1 ;
        RECT 14.065 28.895 14.315 29.905 ;
  LAYER M1 ;
        RECT 13.635 23.015 13.885 26.545 ;
  LAYER M1 ;
        RECT 14.495 23.015 14.745 26.545 ;
  LAYER M1 ;
        RECT 14.925 23.015 15.175 26.545 ;
  LAYER M1 ;
        RECT 14.925 26.795 15.175 27.805 ;
  LAYER M1 ;
        RECT 14.925 28.895 15.175 29.905 ;
  LAYER M1 ;
        RECT 15.355 23.015 15.605 26.545 ;
  LAYER M2 ;
        RECT 14.02 29.26 15.22 29.54 ;
  LAYER M2 ;
        RECT 14.02 22.96 15.22 23.24 ;
  LAYER M2 ;
        RECT 14.02 27.16 15.22 27.44 ;
  LAYER M2 ;
        RECT 13.59 23.38 15.65 23.66 ;
  LAYER M2 ;
        RECT 14.02 37.24 15.22 37.52 ;
  LAYER M2 ;
        RECT 14.02 38.5 15.22 38.78 ;
  LAYER M2 ;
        RECT 18.32 33.04 19.52 33.32 ;
  LAYER M2 ;
        RECT 18.32 42.28 19.52 42.56 ;
  LAYER M2 ;
        RECT 18.76 33.04 19.08 33.32 ;
  LAYER M3 ;
        RECT 18.78 33.18 19.06 42.42 ;
  LAYER M2 ;
        RECT 18.76 42.28 19.08 42.56 ;
  LAYER M2 ;
        RECT 14.46 37.24 14.78 37.52 ;
  LAYER M3 ;
        RECT 14.48 37.38 14.76 38.64 ;
  LAYER M2 ;
        RECT 14.46 38.5 14.78 38.78 ;
  LAYER M3 ;
        RECT 14.48 37.615 14.76 37.985 ;
  LAYER M2 ;
        RECT 14.62 37.66 18.92 37.94 ;
  LAYER M3 ;
        RECT 18.78 37.615 19.06 37.985 ;
  LAYER M2 ;
        RECT 14.46 37.24 14.78 37.52 ;
  LAYER M3 ;
        RECT 14.48 37.22 14.76 37.54 ;
  LAYER M2 ;
        RECT 14.46 38.5 14.78 38.78 ;
  LAYER M3 ;
        RECT 14.48 38.48 14.76 38.8 ;
  LAYER M2 ;
        RECT 14.46 37.24 14.78 37.52 ;
  LAYER M3 ;
        RECT 14.48 37.22 14.76 37.54 ;
  LAYER M2 ;
        RECT 14.46 38.5 14.78 38.78 ;
  LAYER M3 ;
        RECT 14.48 38.48 14.76 38.8 ;
  LAYER M2 ;
        RECT 14.46 37.24 14.78 37.52 ;
  LAYER M3 ;
        RECT 14.48 37.22 14.76 37.54 ;
  LAYER M2 ;
        RECT 14.46 37.66 14.78 37.94 ;
  LAYER M3 ;
        RECT 14.48 37.64 14.76 37.96 ;
  LAYER M2 ;
        RECT 14.46 38.5 14.78 38.78 ;
  LAYER M3 ;
        RECT 14.48 38.48 14.76 38.8 ;
  LAYER M2 ;
        RECT 18.76 37.66 19.08 37.94 ;
  LAYER M3 ;
        RECT 18.78 37.64 19.06 37.96 ;
  LAYER M2 ;
        RECT 14.46 37.24 14.78 37.52 ;
  LAYER M3 ;
        RECT 14.48 37.22 14.76 37.54 ;
  LAYER M2 ;
        RECT 14.46 37.66 14.78 37.94 ;
  LAYER M3 ;
        RECT 14.48 37.64 14.76 37.96 ;
  LAYER M2 ;
        RECT 14.46 38.5 14.78 38.78 ;
  LAYER M3 ;
        RECT 14.48 38.48 14.76 38.8 ;
  LAYER M2 ;
        RECT 18.76 37.66 19.08 37.94 ;
  LAYER M3 ;
        RECT 18.78 37.64 19.06 37.96 ;
  LAYER M2 ;
        RECT 25.2 33.04 26.4 33.32 ;
  LAYER M2 ;
        RECT 25.2 42.28 26.4 42.56 ;
  LAYER M2 ;
        RECT 25.21 33.04 25.53 33.32 ;
  LAYER M3 ;
        RECT 25.23 33.18 25.51 42.42 ;
  LAYER M2 ;
        RECT 25.21 42.28 25.53 42.56 ;
  LAYER M2 ;
        RECT 21.76 37.24 22.96 37.52 ;
  LAYER M2 ;
        RECT 21.76 38.08 22.96 38.36 ;
  LAYER M2 ;
        RECT 22.2 37.24 22.52 37.52 ;
  LAYER M3 ;
        RECT 22.22 37.38 22.5 38.22 ;
  LAYER M2 ;
        RECT 22.2 38.08 22.52 38.36 ;
  LAYER M3 ;
        RECT 25.23 37.615 25.51 37.985 ;
  LAYER M2 ;
        RECT 22.36 37.66 25.37 37.94 ;
  LAYER M3 ;
        RECT 22.22 37.615 22.5 37.985 ;
  LAYER M2 ;
        RECT 22.2 37.66 22.52 37.94 ;
  LAYER M3 ;
        RECT 22.22 37.64 22.5 37.96 ;
  LAYER M2 ;
        RECT 25.21 37.66 25.53 37.94 ;
  LAYER M3 ;
        RECT 25.23 37.64 25.51 37.96 ;
  LAYER M2 ;
        RECT 22.2 37.66 22.52 37.94 ;
  LAYER M3 ;
        RECT 22.22 37.64 22.5 37.96 ;
  LAYER M2 ;
        RECT 25.21 37.66 25.53 37.94 ;
  LAYER M3 ;
        RECT 25.23 37.64 25.51 37.96 ;
  LAYER M2 ;
        RECT 10.58 37.24 11.78 37.52 ;
  LAYER M3 ;
        RECT 14.05 38.06 14.33 42.58 ;
  LAYER M2 ;
        RECT 11.61 37.24 13.33 37.52 ;
  LAYER M3 ;
        RECT 13.19 37.38 13.47 37.8 ;
  LAYER M4 ;
        RECT 13.33 37.4 14.19 38.2 ;
  LAYER M3 ;
        RECT 14.05 37.8 14.33 38.22 ;
  LAYER M2 ;
        RECT 13.17 37.24 13.49 37.52 ;
  LAYER M3 ;
        RECT 13.19 37.22 13.47 37.54 ;
  LAYER M3 ;
        RECT 13.19 37.615 13.47 37.985 ;
  LAYER M4 ;
        RECT 13.165 37.4 13.495 38.2 ;
  LAYER M3 ;
        RECT 14.05 37.615 14.33 37.985 ;
  LAYER M4 ;
        RECT 14.025 37.4 14.355 38.2 ;
  LAYER M2 ;
        RECT 13.17 37.24 13.49 37.52 ;
  LAYER M3 ;
        RECT 13.19 37.22 13.47 37.54 ;
  LAYER M3 ;
        RECT 13.19 37.615 13.47 37.985 ;
  LAYER M4 ;
        RECT 13.165 37.4 13.495 38.2 ;
  LAYER M3 ;
        RECT 14.05 37.615 14.33 37.985 ;
  LAYER M4 ;
        RECT 14.025 37.4 14.355 38.2 ;
  LAYER M2 ;
        RECT 10.15 36.82 12.21 37.1 ;
  LAYER M2 ;
        RECT 9.72 38.08 10.92 38.36 ;
  LAYER M2 ;
        RECT 13.59 36.82 15.65 37.1 ;
  LAYER M2 ;
        RECT 10.16 36.82 10.48 37.1 ;
  LAYER M3 ;
        RECT 10.18 36.96 10.46 38.22 ;
  LAYER M2 ;
        RECT 10.16 38.08 10.48 38.36 ;
  LAYER M2 ;
        RECT 12.04 36.82 13.76 37.1 ;
  LAYER M2 ;
        RECT 10.16 36.82 10.48 37.1 ;
  LAYER M3 ;
        RECT 10.18 36.8 10.46 37.12 ;
  LAYER M2 ;
        RECT 10.16 38.08 10.48 38.36 ;
  LAYER M3 ;
        RECT 10.18 38.06 10.46 38.38 ;
  LAYER M2 ;
        RECT 10.16 36.82 10.48 37.1 ;
  LAYER M3 ;
        RECT 10.18 36.8 10.46 37.12 ;
  LAYER M2 ;
        RECT 10.16 38.08 10.48 38.36 ;
  LAYER M3 ;
        RECT 10.18 38.06 10.46 38.38 ;
  LAYER M2 ;
        RECT 10.16 36.82 10.48 37.1 ;
  LAYER M3 ;
        RECT 10.18 36.8 10.46 37.12 ;
  LAYER M2 ;
        RECT 10.16 38.08 10.48 38.36 ;
  LAYER M3 ;
        RECT 10.18 38.06 10.46 38.38 ;
  LAYER M2 ;
        RECT 10.16 36.82 10.48 37.1 ;
  LAYER M3 ;
        RECT 10.18 36.8 10.46 37.12 ;
  LAYER M2 ;
        RECT 10.16 38.08 10.48 38.36 ;
  LAYER M3 ;
        RECT 10.18 38.06 10.46 38.38 ;
  LAYER M2 ;
        RECT 21.76 33.04 22.96 33.32 ;
  LAYER M2 ;
        RECT 18.32 37.24 19.52 37.52 ;
  LAYER M2 ;
        RECT 18.32 38.08 19.52 38.36 ;
  LAYER M2 ;
        RECT 21.76 42.28 22.96 42.56 ;
  LAYER M2 ;
        RECT 20.64 33.04 21.93 33.32 ;
  LAYER M1 ;
        RECT 20.515 33.18 20.765 37.38 ;
  LAYER M2 ;
        RECT 19.35 37.24 20.64 37.52 ;
  LAYER M2 ;
        RECT 19.19 37.24 19.51 37.52 ;
  LAYER M3 ;
        RECT 19.21 37.38 19.49 38.22 ;
  LAYER M2 ;
        RECT 19.19 38.08 19.51 38.36 ;
  LAYER M1 ;
        RECT 20.515 37.38 20.765 42.42 ;
  LAYER M2 ;
        RECT 20.64 42.28 21.93 42.56 ;
  LAYER M1 ;
        RECT 20.515 33.095 20.765 33.265 ;
  LAYER M2 ;
        RECT 20.47 33.04 20.81 33.32 ;
  LAYER M1 ;
        RECT 20.515 37.295 20.765 37.465 ;
  LAYER M2 ;
        RECT 20.47 37.24 20.81 37.52 ;
  LAYER M1 ;
        RECT 20.515 33.095 20.765 33.265 ;
  LAYER M2 ;
        RECT 20.47 33.04 20.81 33.32 ;
  LAYER M1 ;
        RECT 20.515 37.295 20.765 37.465 ;
  LAYER M2 ;
        RECT 20.47 37.24 20.81 37.52 ;
  LAYER M1 ;
        RECT 20.515 33.095 20.765 33.265 ;
  LAYER M2 ;
        RECT 20.47 33.04 20.81 33.32 ;
  LAYER M1 ;
        RECT 20.515 37.295 20.765 37.465 ;
  LAYER M2 ;
        RECT 20.47 37.24 20.81 37.52 ;
  LAYER M2 ;
        RECT 19.19 37.24 19.51 37.52 ;
  LAYER M3 ;
        RECT 19.21 37.22 19.49 37.54 ;
  LAYER M2 ;
        RECT 19.19 38.08 19.51 38.36 ;
  LAYER M3 ;
        RECT 19.21 38.06 19.49 38.38 ;
  LAYER M1 ;
        RECT 20.515 33.095 20.765 33.265 ;
  LAYER M2 ;
        RECT 20.47 33.04 20.81 33.32 ;
  LAYER M1 ;
        RECT 20.515 37.295 20.765 37.465 ;
  LAYER M2 ;
        RECT 20.47 37.24 20.81 37.52 ;
  LAYER M2 ;
        RECT 19.19 37.24 19.51 37.52 ;
  LAYER M3 ;
        RECT 19.21 37.22 19.49 37.54 ;
  LAYER M2 ;
        RECT 19.19 38.08 19.51 38.36 ;
  LAYER M3 ;
        RECT 19.21 38.06 19.49 38.38 ;
  LAYER M1 ;
        RECT 20.515 33.095 20.765 33.265 ;
  LAYER M2 ;
        RECT 20.47 33.04 20.81 33.32 ;
  LAYER M1 ;
        RECT 20.515 37.295 20.765 37.465 ;
  LAYER M2 ;
        RECT 20.47 37.24 20.81 37.52 ;
  LAYER M1 ;
        RECT 20.515 42.335 20.765 42.505 ;
  LAYER M2 ;
        RECT 20.47 42.28 20.81 42.56 ;
  LAYER M2 ;
        RECT 19.19 37.24 19.51 37.52 ;
  LAYER M3 ;
        RECT 19.21 37.22 19.49 37.54 ;
  LAYER M2 ;
        RECT 19.19 38.08 19.51 38.36 ;
  LAYER M3 ;
        RECT 19.21 38.06 19.49 38.38 ;
  LAYER M1 ;
        RECT 20.515 33.095 20.765 33.265 ;
  LAYER M2 ;
        RECT 20.47 33.04 20.81 33.32 ;
  LAYER M1 ;
        RECT 20.515 37.295 20.765 37.465 ;
  LAYER M2 ;
        RECT 20.47 37.24 20.81 37.52 ;
  LAYER M1 ;
        RECT 20.515 42.335 20.765 42.505 ;
  LAYER M2 ;
        RECT 20.47 42.28 20.81 42.56 ;
  LAYER M2 ;
        RECT 19.19 37.24 19.51 37.52 ;
  LAYER M3 ;
        RECT 19.21 37.22 19.49 37.54 ;
  LAYER M2 ;
        RECT 19.19 38.08 19.51 38.36 ;
  LAYER M3 ;
        RECT 19.21 38.06 19.49 38.38 ;
  LAYER M1 ;
        RECT 19.225 38.135 19.475 41.665 ;
  LAYER M1 ;
        RECT 19.225 41.915 19.475 42.925 ;
  LAYER M1 ;
        RECT 19.225 44.015 19.475 45.025 ;
  LAYER M1 ;
        RECT 19.655 38.135 19.905 41.665 ;
  LAYER M1 ;
        RECT 18.795 38.135 19.045 41.665 ;
  LAYER M1 ;
        RECT 18.365 38.135 18.615 41.665 ;
  LAYER M1 ;
        RECT 18.365 41.915 18.615 42.925 ;
  LAYER M1 ;
        RECT 18.365 44.015 18.615 45.025 ;
  LAYER M1 ;
        RECT 17.935 38.135 18.185 41.665 ;
  LAYER M2 ;
        RECT 17.89 38.5 19.95 38.78 ;
  LAYER M2 ;
        RECT 18.32 44.38 19.52 44.66 ;
  LAYER M2 ;
        RECT 18.32 38.08 19.52 38.36 ;
  LAYER M2 ;
        RECT 18.32 42.28 19.52 42.56 ;
  LAYER M3 ;
        RECT 18.35 38.48 18.63 44.68 ;
  LAYER M1 ;
        RECT 22.665 38.135 22.915 41.665 ;
  LAYER M1 ;
        RECT 22.665 41.915 22.915 42.925 ;
  LAYER M1 ;
        RECT 22.665 44.015 22.915 45.025 ;
  LAYER M1 ;
        RECT 23.095 38.135 23.345 41.665 ;
  LAYER M1 ;
        RECT 22.235 38.135 22.485 41.665 ;
  LAYER M1 ;
        RECT 21.805 38.135 22.055 41.665 ;
  LAYER M1 ;
        RECT 21.805 41.915 22.055 42.925 ;
  LAYER M1 ;
        RECT 21.805 44.015 22.055 45.025 ;
  LAYER M1 ;
        RECT 21.375 38.135 21.625 41.665 ;
  LAYER M2 ;
        RECT 21.33 38.5 23.39 38.78 ;
  LAYER M2 ;
        RECT 21.76 44.38 22.96 44.66 ;
  LAYER M2 ;
        RECT 21.76 38.08 22.96 38.36 ;
  LAYER M2 ;
        RECT 21.76 42.28 22.96 42.56 ;
  LAYER M3 ;
        RECT 21.79 38.48 22.07 44.68 ;
  LAYER M1 ;
        RECT 19.225 33.935 19.475 37.465 ;
  LAYER M1 ;
        RECT 19.225 32.675 19.475 33.685 ;
  LAYER M1 ;
        RECT 19.225 30.575 19.475 31.585 ;
  LAYER M1 ;
        RECT 19.655 33.935 19.905 37.465 ;
  LAYER M1 ;
        RECT 18.795 33.935 19.045 37.465 ;
  LAYER M1 ;
        RECT 18.365 33.935 18.615 37.465 ;
  LAYER M1 ;
        RECT 18.365 32.675 18.615 33.685 ;
  LAYER M1 ;
        RECT 18.365 30.575 18.615 31.585 ;
  LAYER M1 ;
        RECT 17.935 33.935 18.185 37.465 ;
  LAYER M2 ;
        RECT 17.89 36.82 19.95 37.1 ;
  LAYER M2 ;
        RECT 18.32 30.94 19.52 31.22 ;
  LAYER M2 ;
        RECT 18.32 37.24 19.52 37.52 ;
  LAYER M2 ;
        RECT 18.32 33.04 19.52 33.32 ;
  LAYER M3 ;
        RECT 18.35 30.92 18.63 37.12 ;
  LAYER M1 ;
        RECT 22.665 33.935 22.915 37.465 ;
  LAYER M1 ;
        RECT 22.665 32.675 22.915 33.685 ;
  LAYER M1 ;
        RECT 22.665 30.575 22.915 31.585 ;
  LAYER M1 ;
        RECT 23.095 33.935 23.345 37.465 ;
  LAYER M1 ;
        RECT 22.235 33.935 22.485 37.465 ;
  LAYER M1 ;
        RECT 21.805 33.935 22.055 37.465 ;
  LAYER M1 ;
        RECT 21.805 32.675 22.055 33.685 ;
  LAYER M1 ;
        RECT 21.805 30.575 22.055 31.585 ;
  LAYER M1 ;
        RECT 21.375 33.935 21.625 37.465 ;
  LAYER M2 ;
        RECT 21.33 36.82 23.39 37.1 ;
  LAYER M2 ;
        RECT 21.76 30.94 22.96 31.22 ;
  LAYER M2 ;
        RECT 21.76 37.24 22.96 37.52 ;
  LAYER M2 ;
        RECT 21.76 33.04 22.96 33.32 ;
  LAYER M3 ;
        RECT 21.79 30.92 22.07 37.12 ;
  LAYER M1 ;
        RECT 13.205 38.135 13.455 41.665 ;
  LAYER M1 ;
        RECT 13.205 41.915 13.455 42.925 ;
  LAYER M1 ;
        RECT 13.205 44.015 13.455 45.025 ;
  LAYER M1 ;
        RECT 12.775 38.135 13.025 41.665 ;
  LAYER M1 ;
        RECT 13.635 38.135 13.885 41.665 ;
  LAYER M1 ;
        RECT 14.065 38.135 14.315 41.665 ;
  LAYER M1 ;
        RECT 14.065 41.915 14.315 42.925 ;
  LAYER M1 ;
        RECT 14.065 44.015 14.315 45.025 ;
  LAYER M1 ;
        RECT 14.495 38.135 14.745 41.665 ;
  LAYER M1 ;
        RECT 14.925 38.135 15.175 41.665 ;
  LAYER M1 ;
        RECT 14.925 41.915 15.175 42.925 ;
  LAYER M1 ;
        RECT 14.925 44.015 15.175 45.025 ;
  LAYER M1 ;
        RECT 15.355 38.135 15.605 41.665 ;
  LAYER M1 ;
        RECT 15.785 38.135 16.035 41.665 ;
  LAYER M1 ;
        RECT 15.785 41.915 16.035 42.925 ;
  LAYER M1 ;
        RECT 15.785 44.015 16.035 45.025 ;
  LAYER M1 ;
        RECT 16.215 38.135 16.465 41.665 ;
  LAYER M2 ;
        RECT 13.16 38.08 16.08 38.36 ;
  LAYER M2 ;
        RECT 13.16 42.28 16.08 42.56 ;
  LAYER M2 ;
        RECT 12.73 38.92 16.51 39.2 ;
  LAYER M2 ;
        RECT 13.16 44.38 16.08 44.66 ;
  LAYER M3 ;
        RECT 14.05 38.06 14.33 42.58 ;
  LAYER M2 ;
        RECT 14.02 38.5 15.22 38.78 ;
  LAYER M3 ;
        RECT 14.91 38.9 15.19 44.68 ;
  LAYER M1 ;
        RECT 25.245 38.135 25.495 41.665 ;
  LAYER M1 ;
        RECT 25.245 41.915 25.495 42.925 ;
  LAYER M1 ;
        RECT 25.245 44.015 25.495 45.025 ;
  LAYER M1 ;
        RECT 24.815 38.135 25.065 41.665 ;
  LAYER M1 ;
        RECT 25.675 38.135 25.925 41.665 ;
  LAYER M1 ;
        RECT 26.105 38.135 26.355 41.665 ;
  LAYER M1 ;
        RECT 26.105 41.915 26.355 42.925 ;
  LAYER M1 ;
        RECT 26.105 44.015 26.355 45.025 ;
  LAYER M1 ;
        RECT 26.535 38.135 26.785 41.665 ;
  LAYER M2 ;
        RECT 24.77 38.5 26.83 38.78 ;
  LAYER M2 ;
        RECT 25.2 44.38 26.4 44.66 ;
  LAYER M2 ;
        RECT 25.2 38.08 26.4 38.36 ;
  LAYER M2 ;
        RECT 25.2 42.28 26.4 42.56 ;
  LAYER M3 ;
        RECT 26.09 38.48 26.37 44.68 ;
  LAYER M1 ;
        RECT 25.245 33.935 25.495 37.465 ;
  LAYER M1 ;
        RECT 25.245 32.675 25.495 33.685 ;
  LAYER M1 ;
        RECT 25.245 30.575 25.495 31.585 ;
  LAYER M1 ;
        RECT 24.815 33.935 25.065 37.465 ;
  LAYER M1 ;
        RECT 25.675 33.935 25.925 37.465 ;
  LAYER M1 ;
        RECT 26.105 33.935 26.355 37.465 ;
  LAYER M1 ;
        RECT 26.105 32.675 26.355 33.685 ;
  LAYER M1 ;
        RECT 26.105 30.575 26.355 31.585 ;
  LAYER M1 ;
        RECT 26.535 33.935 26.785 37.465 ;
  LAYER M2 ;
        RECT 24.77 36.82 26.83 37.1 ;
  LAYER M2 ;
        RECT 25.2 30.94 26.4 31.22 ;
  LAYER M2 ;
        RECT 25.2 37.24 26.4 37.52 ;
  LAYER M2 ;
        RECT 25.2 33.04 26.4 33.32 ;
  LAYER M3 ;
        RECT 26.09 30.92 26.37 37.12 ;
  LAYER M1 ;
        RECT 9.765 38.135 10.015 41.665 ;
  LAYER M1 ;
        RECT 9.765 41.915 10.015 42.925 ;
  LAYER M1 ;
        RECT 9.765 44.015 10.015 45.025 ;
  LAYER M1 ;
        RECT 9.335 38.135 9.585 41.665 ;
  LAYER M1 ;
        RECT 10.195 38.135 10.445 41.665 ;
  LAYER M1 ;
        RECT 10.625 38.135 10.875 41.665 ;
  LAYER M1 ;
        RECT 10.625 41.915 10.875 42.925 ;
  LAYER M1 ;
        RECT 10.625 44.015 10.875 45.025 ;
  LAYER M1 ;
        RECT 11.055 38.135 11.305 41.665 ;
  LAYER M2 ;
        RECT 9.29 38.5 11.35 38.78 ;
  LAYER M2 ;
        RECT 9.72 44.38 10.92 44.66 ;
  LAYER M2 ;
        RECT 9.72 38.08 10.92 38.36 ;
  LAYER M2 ;
        RECT 9.72 42.28 10.92 42.56 ;
  LAYER M3 ;
        RECT 10.61 38.48 10.89 44.68 ;
  LAYER M1 ;
        RECT 10.625 33.935 10.875 37.465 ;
  LAYER M1 ;
        RECT 10.625 32.675 10.875 33.685 ;
  LAYER M1 ;
        RECT 10.625 30.575 10.875 31.585 ;
  LAYER M1 ;
        RECT 10.195 33.935 10.445 37.465 ;
  LAYER M1 ;
        RECT 11.055 33.935 11.305 37.465 ;
  LAYER M1 ;
        RECT 11.485 33.935 11.735 37.465 ;
  LAYER M1 ;
        RECT 11.485 32.675 11.735 33.685 ;
  LAYER M1 ;
        RECT 11.485 30.575 11.735 31.585 ;
  LAYER M1 ;
        RECT 11.915 33.935 12.165 37.465 ;
  LAYER M2 ;
        RECT 10.58 30.94 11.78 31.22 ;
  LAYER M2 ;
        RECT 10.58 37.24 11.78 37.52 ;
  LAYER M2 ;
        RECT 10.58 33.04 11.78 33.32 ;
  LAYER M2 ;
        RECT 10.15 36.82 12.21 37.1 ;
  LAYER M1 ;
        RECT 14.065 33.935 14.315 37.465 ;
  LAYER M1 ;
        RECT 14.065 32.675 14.315 33.685 ;
  LAYER M1 ;
        RECT 14.065 30.575 14.315 31.585 ;
  LAYER M1 ;
        RECT 13.635 33.935 13.885 37.465 ;
  LAYER M1 ;
        RECT 14.495 33.935 14.745 37.465 ;
  LAYER M1 ;
        RECT 14.925 33.935 15.175 37.465 ;
  LAYER M1 ;
        RECT 14.925 32.675 15.175 33.685 ;
  LAYER M1 ;
        RECT 14.925 30.575 15.175 31.585 ;
  LAYER M1 ;
        RECT 15.355 33.935 15.605 37.465 ;
  LAYER M2 ;
        RECT 14.02 30.94 15.22 31.22 ;
  LAYER M2 ;
        RECT 14.02 37.24 15.22 37.52 ;
  LAYER M2 ;
        RECT 14.02 33.04 15.22 33.32 ;
  LAYER M2 ;
        RECT 13.59 36.82 15.65 37.1 ;
  LAYER M4 ;
        RECT 0.44 24.35 7.74 31.65 ;
  LAYER M4 ;
        RECT 0.44 24.14 0.89 26.66 ;
  LAYER M5 ;
        RECT 7.065 30.67 7.515 33.19 ;
  LAYER M4 ;
        RECT 0.695 32.36 8.335 33.16 ;
  LAYER M4 ;
        RECT 0.695 23.54 8.335 24.34 ;
  LAYER M4 ;
        RECT 0.44 35.69 7.74 42.99 ;
  LAYER M4 ;
        RECT 0.44 35.48 0.89 38 ;
  LAYER M5 ;
        RECT 7.065 42.01 7.515 44.53 ;
  LAYER M4 ;
        RECT 0.695 43.7 8.335 44.5 ;
  LAYER M4 ;
        RECT 0.695 34.88 8.335 35.68 ;
  LAYER M4 ;
        RECT 0.44 1.67 7.74 8.97 ;
  LAYER M4 ;
        RECT 0.44 1.46 0.89 3.98 ;
  LAYER M5 ;
        RECT 7.065 7.99 7.515 10.51 ;
  LAYER M4 ;
        RECT 0.695 9.68 8.335 10.48 ;
  LAYER M4 ;
        RECT 0.695 0.86 8.335 1.66 ;
  LAYER M4 ;
        RECT 0.44 13.01 7.74 20.31 ;
  LAYER M4 ;
        RECT 0.44 12.8 0.89 15.32 ;
  LAYER M5 ;
        RECT 7.065 19.33 7.515 21.85 ;
  LAYER M4 ;
        RECT 0.695 21.02 8.335 21.82 ;
  LAYER M4 ;
        RECT 0.695 12.2 8.335 13 ;
  END 
END TWO_BIT_RES_ADC
