MACRO TWOBIT_DAC
  ORIGIN 0 0 ;
  FOREIGN TWOBIT_DAC 0 0 ;
  SIZE 23.81 BY 23.27 ;
  PIN D0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 19.6 4.9 19.88 ;
      LAYER M2 ;
        RECT 5.42 19.6 6.62 19.88 ;
      LAYER M2 ;
        RECT 4.73 19.6 5.59 19.88 ;
      LAYER M2 ;
        RECT 16.6 19.6 17.8 19.88 ;
      LAYER M2 ;
        RECT 18.32 19.6 19.52 19.88 ;
      LAYER M2 ;
        RECT 17.63 19.6 18.49 19.88 ;
      LAYER M2 ;
        RECT 6.45 19.6 8.17 19.88 ;
      LAYER M1 ;
        RECT 8.045 19.32 8.295 19.74 ;
      LAYER M2 ;
        RECT 8.17 19.18 12.47 19.46 ;
      LAYER M1 ;
        RECT 12.345 19.32 12.595 19.74 ;
      LAYER M2 ;
        RECT 12.47 19.6 16.77 19.88 ;
    END
  END D0
  PIN X2_INP1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.17 6.58 17.37 6.86 ;
      LAYER M2 ;
        RECT 16.6 7.84 17.8 8.12 ;
      LAYER M2 ;
        RECT 16.61 6.58 16.93 6.86 ;
      LAYER M3 ;
        RECT 16.63 6.72 16.91 7.98 ;
      LAYER M2 ;
        RECT 16.61 7.84 16.93 8.12 ;
    END
  END X2_INP1
  PIN X2_INP2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 18.75 6.58 19.95 6.86 ;
      LAYER M2 ;
        RECT 18.32 7.84 19.52 8.12 ;
      LAYER M2 ;
        RECT 18.76 6.58 19.08 6.86 ;
      LAYER M3 ;
        RECT 18.78 6.72 19.06 7.98 ;
      LAYER M2 ;
        RECT 18.76 7.84 19.08 8.12 ;
    END
  END X2_INP2
  PIN X1_INP1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 5.85 6.58 7.05 6.86 ;
      LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
      LAYER M2 ;
        RECT 5.86 6.58 6.18 6.86 ;
      LAYER M3 ;
        RECT 5.88 6.72 6.16 7.98 ;
      LAYER M2 ;
        RECT 5.86 7.84 6.18 8.12 ;
    END
  END X1_INP1
  PIN X1_INP2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
      LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
      LAYER M2 ;
        RECT 4.3 6.58 4.73 6.86 ;
      LAYER M1 ;
        RECT 4.605 6.72 4.855 7.98 ;
      LAYER M2 ;
        RECT 4.57 7.84 4.89 8.12 ;
    END
  END X1_INP2
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.86 19.6 10.06 19.88 ;
      LAYER M2 ;
        RECT 10.58 19.6 11.78 19.88 ;
      LAYER M2 ;
        RECT 9.89 19.6 10.75 19.88 ;
    END
  END D1
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
      LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
      LAYER M2 ;
        RECT 10.58 7 11.78 7.28 ;
      LAYER M2 ;
        RECT 11.01 8.26 12.21 8.54 ;
      LAYER M2 ;
        RECT 9.3 7 9.62 7.28 ;
      LAYER M3 ;
        RECT 9.32 7.14 9.6 8.4 ;
      LAYER M2 ;
        RECT 9.3 8.26 9.62 8.54 ;
      LAYER M2 ;
        RECT 9.89 7 10.75 7.28 ;
      LAYER M2 ;
        RECT 9.46 8.26 11.18 8.54 ;
    END
  END OUT
  OBS 
  LAYER M2 ;
        RECT 11.01 6.58 12.21 6.86 ;
  LAYER M2 ;
        RECT 10.58 7.84 11.78 8.12 ;
  LAYER M2 ;
        RECT 11.02 6.58 11.34 6.86 ;
  LAYER M3 ;
        RECT 11.04 6.72 11.32 7.98 ;
  LAYER M2 ;
        RECT 11.02 7.84 11.34 8.12 ;
  LAYER M2 ;
        RECT 16.6 7 17.8 7.28 ;
  LAYER M2 ;
        RECT 16.17 8.26 17.37 8.54 ;
  LAYER M2 ;
        RECT 18.32 7 19.52 7.28 ;
  LAYER M2 ;
        RECT 18.75 8.26 19.95 8.54 ;
  LAYER M2 ;
        RECT 17.04 7 17.36 7.28 ;
  LAYER M3 ;
        RECT 17.06 7.14 17.34 8.4 ;
  LAYER M2 ;
        RECT 17.04 8.26 17.36 8.54 ;
  LAYER M2 ;
        RECT 17.63 7 18.49 7.28 ;
  LAYER M2 ;
        RECT 17.2 8.26 18.92 8.54 ;
  LAYER M2 ;
        RECT 11.61 7.84 15.91 8.12 ;
  LAYER M3 ;
        RECT 15.77 7.98 16.05 8.4 ;
  LAYER M2 ;
        RECT 15.91 8.26 16.34 8.54 ;
  LAYER M2 ;
        RECT 15.75 7.84 16.07 8.12 ;
  LAYER M3 ;
        RECT 15.77 7.82 16.05 8.14 ;
  LAYER M2 ;
        RECT 15.75 8.26 16.07 8.54 ;
  LAYER M3 ;
        RECT 15.77 8.24 16.05 8.56 ;
  LAYER M2 ;
        RECT 15.75 7.84 16.07 8.12 ;
  LAYER M3 ;
        RECT 15.77 7.82 16.05 8.14 ;
  LAYER M2 ;
        RECT 15.75 8.26 16.07 8.54 ;
  LAYER M3 ;
        RECT 15.77 8.24 16.05 8.56 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 4.14 7 4.46 7.28 ;
  LAYER M3 ;
        RECT 4.16 7.14 4.44 8.4 ;
  LAYER M2 ;
        RECT 4.14 8.26 4.46 8.54 ;
  LAYER M2 ;
        RECT 4.73 7 5.59 7.28 ;
  LAYER M2 ;
        RECT 4.3 8.26 6.02 8.54 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8.86 7.84 10.06 8.12 ;
  LAYER M2 ;
        RECT 8.87 6.58 9.19 6.86 ;
  LAYER M3 ;
        RECT 8.89 6.72 9.17 7.98 ;
  LAYER M2 ;
        RECT 8.87 7.84 9.19 8.12 ;
  LAYER M2 ;
        RECT 6.88 8.26 7.74 8.54 ;
  LAYER M3 ;
        RECT 7.6 7.98 7.88 8.4 ;
  LAYER M2 ;
        RECT 7.74 7.84 9.03 8.12 ;
  LAYER M2 ;
        RECT 7.58 7.84 7.9 8.12 ;
  LAYER M3 ;
        RECT 7.6 7.82 7.88 8.14 ;
  LAYER M2 ;
        RECT 7.58 8.26 7.9 8.54 ;
  LAYER M3 ;
        RECT 7.6 8.24 7.88 8.56 ;
  LAYER M2 ;
        RECT 7.58 7.84 7.9 8.12 ;
  LAYER M3 ;
        RECT 7.6 7.82 7.88 8.14 ;
  LAYER M2 ;
        RECT 7.58 8.26 7.9 8.54 ;
  LAYER M3 ;
        RECT 7.6 8.24 7.88 8.56 ;
  LAYER M2 ;
        RECT 16.6 2.8 17.8 3.08 ;
  LAYER M2 ;
        RECT 18.32 2.8 19.52 3.08 ;
  LAYER M2 ;
        RECT 20.9 6.16 22.1 6.44 ;
  LAYER M2 ;
        RECT 20.9 15.4 22.1 15.68 ;
  LAYER M2 ;
        RECT 18.32 15.4 19.52 15.68 ;
  LAYER M2 ;
        RECT 16.6 15.4 17.8 15.68 ;
  LAYER M2 ;
        RECT 17.63 2.8 18.49 3.08 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.94 19.49 6.3 ;
  LAYER M2 ;
        RECT 19.35 6.16 21.07 6.44 ;
  LAYER M2 ;
        RECT 20.91 6.16 21.23 6.44 ;
  LAYER M1 ;
        RECT 20.945 6.3 21.195 15.54 ;
  LAYER M2 ;
        RECT 20.91 15.4 21.23 15.68 ;
  LAYER M2 ;
        RECT 19.35 15.4 21.07 15.68 ;
  LAYER M2 ;
        RECT 17.63 15.4 18.49 15.68 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.78 19.49 3.1 ;
  LAYER M2 ;
        RECT 19.19 6.16 19.51 6.44 ;
  LAYER M3 ;
        RECT 19.21 6.14 19.49 6.46 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.78 19.49 3.1 ;
  LAYER M2 ;
        RECT 19.19 6.16 19.51 6.44 ;
  LAYER M3 ;
        RECT 19.21 6.14 19.49 6.46 ;
  LAYER M1 ;
        RECT 20.945 6.215 21.195 6.385 ;
  LAYER M2 ;
        RECT 20.9 6.16 21.24 6.44 ;
  LAYER M1 ;
        RECT 20.945 15.455 21.195 15.625 ;
  LAYER M2 ;
        RECT 20.9 15.4 21.24 15.68 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.78 19.49 3.1 ;
  LAYER M2 ;
        RECT 19.19 6.16 19.51 6.44 ;
  LAYER M3 ;
        RECT 19.21 6.14 19.49 6.46 ;
  LAYER M1 ;
        RECT 20.945 6.215 21.195 6.385 ;
  LAYER M2 ;
        RECT 20.9 6.16 21.24 6.44 ;
  LAYER M1 ;
        RECT 20.945 15.455 21.195 15.625 ;
  LAYER M2 ;
        RECT 20.9 15.4 21.24 15.68 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.78 19.49 3.1 ;
  LAYER M2 ;
        RECT 19.19 6.16 19.51 6.44 ;
  LAYER M3 ;
        RECT 19.21 6.14 19.49 6.46 ;
  LAYER M1 ;
        RECT 20.945 6.215 21.195 6.385 ;
  LAYER M2 ;
        RECT 20.9 6.16 21.24 6.44 ;
  LAYER M1 ;
        RECT 20.945 15.455 21.195 15.625 ;
  LAYER M2 ;
        RECT 20.9 15.4 21.24 15.68 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.78 19.49 3.1 ;
  LAYER M2 ;
        RECT 19.19 6.16 19.51 6.44 ;
  LAYER M3 ;
        RECT 19.21 6.14 19.49 6.46 ;
  LAYER M1 ;
        RECT 20.945 6.215 21.195 6.385 ;
  LAYER M2 ;
        RECT 20.9 6.16 21.24 6.44 ;
  LAYER M1 ;
        RECT 20.945 15.455 21.195 15.625 ;
  LAYER M2 ;
        RECT 20.9 15.4 21.24 15.68 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.78 19.49 3.1 ;
  LAYER M2 ;
        RECT 19.19 6.16 19.51 6.44 ;
  LAYER M3 ;
        RECT 19.21 6.14 19.49 6.46 ;
  LAYER M1 ;
        RECT 20.945 6.215 21.195 6.385 ;
  LAYER M2 ;
        RECT 20.9 6.16 21.24 6.44 ;
  LAYER M1 ;
        RECT 20.945 15.455 21.195 15.625 ;
  LAYER M2 ;
        RECT 20.9 15.4 21.24 15.68 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.78 19.49 3.1 ;
  LAYER M2 ;
        RECT 19.19 6.16 19.51 6.44 ;
  LAYER M3 ;
        RECT 19.21 6.14 19.49 6.46 ;
  LAYER M1 ;
        RECT 20.945 6.215 21.195 6.385 ;
  LAYER M2 ;
        RECT 20.9 6.16 21.24 6.44 ;
  LAYER M1 ;
        RECT 20.945 15.455 21.195 15.625 ;
  LAYER M2 ;
        RECT 20.9 15.4 21.24 15.68 ;
  LAYER M2 ;
        RECT 19.19 2.8 19.51 3.08 ;
  LAYER M3 ;
        RECT 19.21 2.78 19.49 3.1 ;
  LAYER M2 ;
        RECT 19.19 6.16 19.51 6.44 ;
  LAYER M3 ;
        RECT 19.21 6.14 19.49 6.46 ;
  LAYER M2 ;
        RECT 16.6 12.04 17.8 12.32 ;
  LAYER M2 ;
        RECT 18.32 12.04 19.52 12.32 ;
  LAYER M2 ;
        RECT 20.9 11.2 22.1 11.48 ;
  LAYER M2 ;
        RECT 20.9 10.36 22.1 10.64 ;
  LAYER M2 ;
        RECT 17.63 12.04 18.49 12.32 ;
  LAYER M2 ;
        RECT 19.35 12.04 19.78 12.32 ;
  LAYER M3 ;
        RECT 19.64 11.34 19.92 12.18 ;
  LAYER M2 ;
        RECT 19.78 11.2 21.07 11.48 ;
  LAYER M2 ;
        RECT 20.91 11.2 21.23 11.48 ;
  LAYER M3 ;
        RECT 20.93 10.5 21.21 11.34 ;
  LAYER M2 ;
        RECT 20.91 10.36 21.23 10.64 ;
  LAYER M2 ;
        RECT 19.62 11.2 19.94 11.48 ;
  LAYER M3 ;
        RECT 19.64 11.18 19.92 11.5 ;
  LAYER M2 ;
        RECT 19.62 12.04 19.94 12.32 ;
  LAYER M3 ;
        RECT 19.64 12.02 19.92 12.34 ;
  LAYER M2 ;
        RECT 19.62 11.2 19.94 11.48 ;
  LAYER M3 ;
        RECT 19.64 11.18 19.92 11.5 ;
  LAYER M2 ;
        RECT 19.62 12.04 19.94 12.32 ;
  LAYER M3 ;
        RECT 19.64 12.02 19.92 12.34 ;
  LAYER M2 ;
        RECT 19.62 11.2 19.94 11.48 ;
  LAYER M3 ;
        RECT 19.64 11.18 19.92 11.5 ;
  LAYER M2 ;
        RECT 19.62 12.04 19.94 12.32 ;
  LAYER M3 ;
        RECT 19.64 12.02 19.92 12.34 ;
  LAYER M2 ;
        RECT 20.91 10.36 21.23 10.64 ;
  LAYER M3 ;
        RECT 20.93 10.34 21.21 10.66 ;
  LAYER M2 ;
        RECT 20.91 11.2 21.23 11.48 ;
  LAYER M3 ;
        RECT 20.93 11.18 21.21 11.5 ;
  LAYER M2 ;
        RECT 19.62 11.2 19.94 11.48 ;
  LAYER M3 ;
        RECT 19.64 11.18 19.92 11.5 ;
  LAYER M2 ;
        RECT 19.62 12.04 19.94 12.32 ;
  LAYER M3 ;
        RECT 19.64 12.02 19.92 12.34 ;
  LAYER M2 ;
        RECT 20.91 10.36 21.23 10.64 ;
  LAYER M3 ;
        RECT 20.93 10.34 21.21 10.66 ;
  LAYER M2 ;
        RECT 20.91 11.2 21.23 11.48 ;
  LAYER M3 ;
        RECT 20.93 11.18 21.21 11.5 ;
  LAYER M1 ;
        RECT 19.225 15.455 19.475 18.985 ;
  LAYER M1 ;
        RECT 19.225 19.235 19.475 20.245 ;
  LAYER M1 ;
        RECT 19.225 21.335 19.475 22.345 ;
  LAYER M1 ;
        RECT 18.795 15.455 19.045 18.985 ;
  LAYER M1 ;
        RECT 19.655 15.455 19.905 18.985 ;
  LAYER M2 ;
        RECT 18.75 21.7 19.95 21.98 ;
  LAYER M2 ;
        RECT 18.75 15.82 19.95 16.1 ;
  LAYER M2 ;
        RECT 18.32 15.4 19.52 15.68 ;
  LAYER M2 ;
        RECT 18.32 19.6 19.52 19.88 ;
  LAYER M3 ;
        RECT 19.64 15.8 19.92 22 ;
  LAYER M1 ;
        RECT 21.805 11.255 22.055 14.785 ;
  LAYER M1 ;
        RECT 21.805 15.035 22.055 16.045 ;
  LAYER M1 ;
        RECT 21.805 17.135 22.055 18.145 ;
  LAYER M1 ;
        RECT 21.375 11.255 21.625 14.785 ;
  LAYER M1 ;
        RECT 22.235 11.255 22.485 14.785 ;
  LAYER M2 ;
        RECT 21.33 17.5 22.53 17.78 ;
  LAYER M2 ;
        RECT 21.33 11.62 22.53 11.9 ;
  LAYER M2 ;
        RECT 20.9 11.2 22.1 11.48 ;
  LAYER M2 ;
        RECT 20.9 15.4 22.1 15.68 ;
  LAYER M3 ;
        RECT 22.22 11.6 22.5 17.8 ;
  LAYER M1 ;
        RECT 16.645 15.455 16.895 18.985 ;
  LAYER M1 ;
        RECT 16.645 19.235 16.895 20.245 ;
  LAYER M1 ;
        RECT 16.645 21.335 16.895 22.345 ;
  LAYER M1 ;
        RECT 17.075 15.455 17.325 18.985 ;
  LAYER M1 ;
        RECT 16.215 15.455 16.465 18.985 ;
  LAYER M2 ;
        RECT 16.17 21.7 17.37 21.98 ;
  LAYER M2 ;
        RECT 16.17 15.82 17.37 16.1 ;
  LAYER M2 ;
        RECT 16.6 15.4 17.8 15.68 ;
  LAYER M2 ;
        RECT 16.6 19.6 17.8 19.88 ;
  LAYER M3 ;
        RECT 16.2 15.8 16.48 22 ;
  LAYER M1 ;
        RECT 21.805 7.055 22.055 10.585 ;
  LAYER M1 ;
        RECT 21.805 5.795 22.055 6.805 ;
  LAYER M1 ;
        RECT 21.805 3.695 22.055 4.705 ;
  LAYER M1 ;
        RECT 21.375 7.055 21.625 10.585 ;
  LAYER M1 ;
        RECT 22.235 7.055 22.485 10.585 ;
  LAYER M2 ;
        RECT 21.33 4.06 22.53 4.34 ;
  LAYER M2 ;
        RECT 21.33 9.94 22.53 10.22 ;
  LAYER M2 ;
        RECT 20.9 10.36 22.1 10.64 ;
  LAYER M2 ;
        RECT 20.9 6.16 22.1 6.44 ;
  LAYER M3 ;
        RECT 22.22 4.04 22.5 10.24 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 12.685 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 14.785 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M2 ;
        RECT 16.6 14.14 17.8 14.42 ;
  LAYER M2 ;
        RECT 16.6 7.84 17.8 8.12 ;
  LAYER M2 ;
        RECT 16.6 12.04 17.8 12.32 ;
  LAYER M2 ;
        RECT 16.17 8.26 17.37 8.54 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M2 ;
        RECT 18.32 0.7 19.52 0.98 ;
  LAYER M2 ;
        RECT 18.32 7 19.52 7.28 ;
  LAYER M2 ;
        RECT 18.32 2.8 19.52 3.08 ;
  LAYER M2 ;
        RECT 18.75 6.58 19.95 6.86 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 11.425 ;
  LAYER M1 ;
        RECT 19.225 11.675 19.475 12.685 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 14.785 ;
  LAYER M1 ;
        RECT 18.795 7.895 19.045 11.425 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M2 ;
        RECT 18.32 14.14 19.52 14.42 ;
  LAYER M2 ;
        RECT 18.32 7.84 19.52 8.12 ;
  LAYER M2 ;
        RECT 18.32 12.04 19.52 12.32 ;
  LAYER M2 ;
        RECT 18.75 8.26 19.95 8.54 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M2 ;
        RECT 16.6 0.7 17.8 0.98 ;
  LAYER M2 ;
        RECT 16.6 7 17.8 7.28 ;
  LAYER M2 ;
        RECT 16.6 2.8 17.8 3.08 ;
  LAYER M2 ;
        RECT 16.17 6.58 17.37 6.86 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
  LAYER M2 ;
        RECT 1.12 6.16 2.32 6.44 ;
  LAYER M2 ;
        RECT 1.12 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 3.7 15.4 4.9 15.68 ;
  LAYER M2 ;
        RECT 5.42 15.4 6.62 15.68 ;
  LAYER M2 ;
        RECT 4.73 2.8 5.59 3.08 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.94 4.01 6.3 ;
  LAYER M2 ;
        RECT 2.15 6.16 3.87 6.44 ;
  LAYER M2 ;
        RECT 1.99 6.16 2.31 6.44 ;
  LAYER M1 ;
        RECT 2.025 6.3 2.275 15.54 ;
  LAYER M2 ;
        RECT 1.99 15.4 2.31 15.68 ;
  LAYER M2 ;
        RECT 2.15 15.4 3.87 15.68 ;
  LAYER M2 ;
        RECT 4.73 15.4 5.59 15.68 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 3.1 ;
  LAYER M2 ;
        RECT 3.71 6.16 4.03 6.44 ;
  LAYER M3 ;
        RECT 3.73 6.14 4.01 6.46 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 3.1 ;
  LAYER M2 ;
        RECT 3.71 6.16 4.03 6.44 ;
  LAYER M3 ;
        RECT 3.73 6.14 4.01 6.46 ;
  LAYER M1 ;
        RECT 2.025 6.215 2.275 6.385 ;
  LAYER M2 ;
        RECT 1.98 6.16 2.32 6.44 ;
  LAYER M1 ;
        RECT 2.025 15.455 2.275 15.625 ;
  LAYER M2 ;
        RECT 1.98 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 3.1 ;
  LAYER M2 ;
        RECT 3.71 6.16 4.03 6.44 ;
  LAYER M3 ;
        RECT 3.73 6.14 4.01 6.46 ;
  LAYER M1 ;
        RECT 2.025 6.215 2.275 6.385 ;
  LAYER M2 ;
        RECT 1.98 6.16 2.32 6.44 ;
  LAYER M1 ;
        RECT 2.025 15.455 2.275 15.625 ;
  LAYER M2 ;
        RECT 1.98 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 3.1 ;
  LAYER M2 ;
        RECT 3.71 6.16 4.03 6.44 ;
  LAYER M3 ;
        RECT 3.73 6.14 4.01 6.46 ;
  LAYER M1 ;
        RECT 2.025 6.215 2.275 6.385 ;
  LAYER M2 ;
        RECT 1.98 6.16 2.32 6.44 ;
  LAYER M1 ;
        RECT 2.025 15.455 2.275 15.625 ;
  LAYER M2 ;
        RECT 1.98 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 3.1 ;
  LAYER M2 ;
        RECT 3.71 6.16 4.03 6.44 ;
  LAYER M3 ;
        RECT 3.73 6.14 4.01 6.46 ;
  LAYER M1 ;
        RECT 2.025 6.215 2.275 6.385 ;
  LAYER M2 ;
        RECT 1.98 6.16 2.32 6.44 ;
  LAYER M1 ;
        RECT 2.025 15.455 2.275 15.625 ;
  LAYER M2 ;
        RECT 1.98 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 3.1 ;
  LAYER M2 ;
        RECT 3.71 6.16 4.03 6.44 ;
  LAYER M3 ;
        RECT 3.73 6.14 4.01 6.46 ;
  LAYER M1 ;
        RECT 2.025 6.215 2.275 6.385 ;
  LAYER M2 ;
        RECT 1.98 6.16 2.32 6.44 ;
  LAYER M1 ;
        RECT 2.025 15.455 2.275 15.625 ;
  LAYER M2 ;
        RECT 1.98 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 3.1 ;
  LAYER M2 ;
        RECT 3.71 6.16 4.03 6.44 ;
  LAYER M3 ;
        RECT 3.73 6.14 4.01 6.46 ;
  LAYER M1 ;
        RECT 2.025 6.215 2.275 6.385 ;
  LAYER M2 ;
        RECT 1.98 6.16 2.32 6.44 ;
  LAYER M1 ;
        RECT 2.025 15.455 2.275 15.625 ;
  LAYER M2 ;
        RECT 1.98 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
  LAYER M3 ;
        RECT 3.73 2.78 4.01 3.1 ;
  LAYER M2 ;
        RECT 3.71 6.16 4.03 6.44 ;
  LAYER M3 ;
        RECT 3.73 6.14 4.01 6.46 ;
  LAYER M2 ;
        RECT 1.12 10.36 2.32 10.64 ;
  LAYER M2 ;
        RECT 1.12 11.2 2.32 11.48 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.5 2.29 11.34 ;
  LAYER M2 ;
        RECT 1.99 11.2 2.31 11.48 ;
  LAYER M3 ;
        RECT 2.01 11.34 2.29 12.18 ;
  LAYER M2 ;
        RECT 2.15 12.04 3.87 12.32 ;
  LAYER M2 ;
        RECT 4.73 12.04 5.59 12.32 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 11.2 2.31 11.48 ;
  LAYER M3 ;
        RECT 2.01 11.18 2.29 11.5 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 11.2 2.31 11.48 ;
  LAYER M3 ;
        RECT 2.01 11.18 2.29 11.5 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 11.2 2.31 11.48 ;
  LAYER M3 ;
        RECT 2.01 11.18 2.29 11.5 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 11.2 2.31 11.48 ;
  LAYER M3 ;
        RECT 2.01 11.18 2.29 11.5 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 11.2 2.31 11.48 ;
  LAYER M3 ;
        RECT 2.01 11.18 2.29 11.5 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 11.2 2.31 11.48 ;
  LAYER M3 ;
        RECT 2.01 11.18 2.29 11.5 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 18.985 ;
  LAYER M1 ;
        RECT 3.745 19.235 3.995 20.245 ;
  LAYER M1 ;
        RECT 3.745 21.335 3.995 22.345 ;
  LAYER M1 ;
        RECT 4.175 15.455 4.425 18.985 ;
  LAYER M1 ;
        RECT 3.315 15.455 3.565 18.985 ;
  LAYER M2 ;
        RECT 3.27 21.7 4.47 21.98 ;
  LAYER M2 ;
        RECT 3.27 15.82 4.47 16.1 ;
  LAYER M2 ;
        RECT 3.7 15.4 4.9 15.68 ;
  LAYER M2 ;
        RECT 3.7 19.6 4.9 19.88 ;
  LAYER M3 ;
        RECT 3.3 15.8 3.58 22 ;
  LAYER M1 ;
        RECT 1.165 11.255 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.165 15.035 1.415 16.045 ;
  LAYER M1 ;
        RECT 1.165 17.135 1.415 18.145 ;
  LAYER M1 ;
        RECT 1.595 11.255 1.845 14.785 ;
  LAYER M1 ;
        RECT 0.735 11.255 0.985 14.785 ;
  LAYER M2 ;
        RECT 0.69 17.5 1.89 17.78 ;
  LAYER M2 ;
        RECT 0.69 11.62 1.89 11.9 ;
  LAYER M2 ;
        RECT 1.12 11.2 2.32 11.48 ;
  LAYER M2 ;
        RECT 1.12 15.4 2.32 15.68 ;
  LAYER M3 ;
        RECT 0.72 11.6 1 17.8 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 18.985 ;
  LAYER M1 ;
        RECT 6.325 19.235 6.575 20.245 ;
  LAYER M1 ;
        RECT 6.325 21.335 6.575 22.345 ;
  LAYER M1 ;
        RECT 5.895 15.455 6.145 18.985 ;
  LAYER M1 ;
        RECT 6.755 15.455 7.005 18.985 ;
  LAYER M2 ;
        RECT 5.85 21.7 7.05 21.98 ;
  LAYER M2 ;
        RECT 5.85 15.82 7.05 16.1 ;
  LAYER M2 ;
        RECT 5.42 15.4 6.62 15.68 ;
  LAYER M2 ;
        RECT 5.42 19.6 6.62 19.88 ;
  LAYER M3 ;
        RECT 6.74 15.8 7.02 22 ;
  LAYER M1 ;
        RECT 1.165 7.055 1.415 10.585 ;
  LAYER M1 ;
        RECT 1.165 5.795 1.415 6.805 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 4.705 ;
  LAYER M1 ;
        RECT 1.595 7.055 1.845 10.585 ;
  LAYER M1 ;
        RECT 0.735 7.055 0.985 10.585 ;
  LAYER M2 ;
        RECT 0.69 4.06 1.89 4.34 ;
  LAYER M2 ;
        RECT 0.69 9.94 1.89 10.22 ;
  LAYER M2 ;
        RECT 1.12 10.36 2.32 10.64 ;
  LAYER M2 ;
        RECT 1.12 6.16 2.32 6.44 ;
  LAYER M3 ;
        RECT 0.72 4.04 1 10.24 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M2 ;
        RECT 5.42 14.14 6.62 14.42 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.7 0.7 4.9 0.98 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M2 ;
        RECT 3.7 14.14 4.9 14.42 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 5.42 0.7 6.62 0.98 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
  LAYER M2 ;
        RECT 5.85 6.58 7.05 6.86 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M2 ;
        RECT 10.58 2.8 11.78 3.08 ;
  LAYER M2 ;
        RECT 13.16 6.16 14.36 6.44 ;
  LAYER M2 ;
        RECT 13.16 15.4 14.36 15.68 ;
  LAYER M2 ;
        RECT 10.58 15.4 11.78 15.68 ;
  LAYER M2 ;
        RECT 8.86 15.4 10.06 15.68 ;
  LAYER M2 ;
        RECT 9.89 2.8 10.75 3.08 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.94 11.75 6.3 ;
  LAYER M2 ;
        RECT 11.61 6.16 13.33 6.44 ;
  LAYER M2 ;
        RECT 13.17 6.16 13.49 6.44 ;
  LAYER M1 ;
        RECT 13.205 6.3 13.455 15.54 ;
  LAYER M2 ;
        RECT 13.17 15.4 13.49 15.68 ;
  LAYER M2 ;
        RECT 11.61 15.4 13.33 15.68 ;
  LAYER M2 ;
        RECT 9.89 15.4 10.75 15.68 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 3.1 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 3.1 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M1 ;
        RECT 13.205 6.215 13.455 6.385 ;
  LAYER M2 ;
        RECT 13.16 6.16 13.5 6.44 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 15.625 ;
  LAYER M2 ;
        RECT 13.16 15.4 13.5 15.68 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 3.1 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M1 ;
        RECT 13.205 6.215 13.455 6.385 ;
  LAYER M2 ;
        RECT 13.16 6.16 13.5 6.44 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 15.625 ;
  LAYER M2 ;
        RECT 13.16 15.4 13.5 15.68 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 3.1 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M1 ;
        RECT 13.205 6.215 13.455 6.385 ;
  LAYER M2 ;
        RECT 13.16 6.16 13.5 6.44 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 15.625 ;
  LAYER M2 ;
        RECT 13.16 15.4 13.5 15.68 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 3.1 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M1 ;
        RECT 13.205 6.215 13.455 6.385 ;
  LAYER M2 ;
        RECT 13.16 6.16 13.5 6.44 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 15.625 ;
  LAYER M2 ;
        RECT 13.16 15.4 13.5 15.68 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 3.1 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M1 ;
        RECT 13.205 6.215 13.455 6.385 ;
  LAYER M2 ;
        RECT 13.16 6.16 13.5 6.44 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 15.625 ;
  LAYER M2 ;
        RECT 13.16 15.4 13.5 15.68 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 3.1 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M1 ;
        RECT 13.205 6.215 13.455 6.385 ;
  LAYER M2 ;
        RECT 13.16 6.16 13.5 6.44 ;
  LAYER M1 ;
        RECT 13.205 15.455 13.455 15.625 ;
  LAYER M2 ;
        RECT 13.16 15.4 13.5 15.68 ;
  LAYER M2 ;
        RECT 11.45 2.8 11.77 3.08 ;
  LAYER M3 ;
        RECT 11.47 2.78 11.75 3.1 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.06 12.32 ;
  LAYER M2 ;
        RECT 10.58 12.04 11.78 12.32 ;
  LAYER M2 ;
        RECT 13.16 11.2 14.36 11.48 ;
  LAYER M2 ;
        RECT 13.16 10.36 14.36 10.64 ;
  LAYER M2 ;
        RECT 9.89 12.04 10.75 12.32 ;
  LAYER M2 ;
        RECT 11.61 12.04 12.04 12.32 ;
  LAYER M3 ;
        RECT 11.9 11.34 12.18 12.18 ;
  LAYER M2 ;
        RECT 12.04 11.2 13.33 11.48 ;
  LAYER M2 ;
        RECT 13.17 11.2 13.49 11.48 ;
  LAYER M3 ;
        RECT 13.19 10.5 13.47 11.34 ;
  LAYER M2 ;
        RECT 13.17 10.36 13.49 10.64 ;
  LAYER M2 ;
        RECT 11.88 11.2 12.2 11.48 ;
  LAYER M3 ;
        RECT 11.9 11.18 12.18 11.5 ;
  LAYER M2 ;
        RECT 11.88 12.04 12.2 12.32 ;
  LAYER M3 ;
        RECT 11.9 12.02 12.18 12.34 ;
  LAYER M2 ;
        RECT 11.88 11.2 12.2 11.48 ;
  LAYER M3 ;
        RECT 11.9 11.18 12.18 11.5 ;
  LAYER M2 ;
        RECT 11.88 12.04 12.2 12.32 ;
  LAYER M3 ;
        RECT 11.9 12.02 12.18 12.34 ;
  LAYER M2 ;
        RECT 11.88 11.2 12.2 11.48 ;
  LAYER M3 ;
        RECT 11.9 11.18 12.18 11.5 ;
  LAYER M2 ;
        RECT 11.88 12.04 12.2 12.32 ;
  LAYER M3 ;
        RECT 11.9 12.02 12.18 12.34 ;
  LAYER M2 ;
        RECT 13.17 10.36 13.49 10.64 ;
  LAYER M3 ;
        RECT 13.19 10.34 13.47 10.66 ;
  LAYER M2 ;
        RECT 13.17 11.2 13.49 11.48 ;
  LAYER M3 ;
        RECT 13.19 11.18 13.47 11.5 ;
  LAYER M2 ;
        RECT 11.88 11.2 12.2 11.48 ;
  LAYER M3 ;
        RECT 11.9 11.18 12.18 11.5 ;
  LAYER M2 ;
        RECT 11.88 12.04 12.2 12.32 ;
  LAYER M3 ;
        RECT 11.9 12.02 12.18 12.34 ;
  LAYER M2 ;
        RECT 13.17 10.36 13.49 10.64 ;
  LAYER M3 ;
        RECT 13.19 10.34 13.47 10.66 ;
  LAYER M2 ;
        RECT 13.17 11.2 13.49 11.48 ;
  LAYER M3 ;
        RECT 13.19 11.18 13.47 11.5 ;
  LAYER M1 ;
        RECT 11.485 15.455 11.735 18.985 ;
  LAYER M1 ;
        RECT 11.485 19.235 11.735 20.245 ;
  LAYER M1 ;
        RECT 11.485 21.335 11.735 22.345 ;
  LAYER M1 ;
        RECT 11.055 15.455 11.305 18.985 ;
  LAYER M1 ;
        RECT 11.915 15.455 12.165 18.985 ;
  LAYER M2 ;
        RECT 11.01 21.7 12.21 21.98 ;
  LAYER M2 ;
        RECT 11.01 15.82 12.21 16.1 ;
  LAYER M2 ;
        RECT 10.58 15.4 11.78 15.68 ;
  LAYER M2 ;
        RECT 10.58 19.6 11.78 19.88 ;
  LAYER M3 ;
        RECT 11.9 15.8 12.18 22 ;
  LAYER M1 ;
        RECT 14.065 11.255 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.065 15.035 14.315 16.045 ;
  LAYER M1 ;
        RECT 14.065 17.135 14.315 18.145 ;
  LAYER M1 ;
        RECT 13.635 11.255 13.885 14.785 ;
  LAYER M1 ;
        RECT 14.495 11.255 14.745 14.785 ;
  LAYER M2 ;
        RECT 13.59 17.5 14.79 17.78 ;
  LAYER M2 ;
        RECT 13.59 11.62 14.79 11.9 ;
  LAYER M2 ;
        RECT 13.16 11.2 14.36 11.48 ;
  LAYER M2 ;
        RECT 13.16 15.4 14.36 15.68 ;
  LAYER M3 ;
        RECT 14.48 11.6 14.76 17.8 ;
  LAYER M1 ;
        RECT 8.905 15.455 9.155 18.985 ;
  LAYER M1 ;
        RECT 8.905 19.235 9.155 20.245 ;
  LAYER M1 ;
        RECT 8.905 21.335 9.155 22.345 ;
  LAYER M1 ;
        RECT 9.335 15.455 9.585 18.985 ;
  LAYER M1 ;
        RECT 8.475 15.455 8.725 18.985 ;
  LAYER M2 ;
        RECT 8.43 21.7 9.63 21.98 ;
  LAYER M2 ;
        RECT 8.43 15.82 9.63 16.1 ;
  LAYER M2 ;
        RECT 8.86 15.4 10.06 15.68 ;
  LAYER M2 ;
        RECT 8.86 19.6 10.06 19.88 ;
  LAYER M3 ;
        RECT 8.46 15.8 8.74 22 ;
  LAYER M1 ;
        RECT 14.065 7.055 14.315 10.585 ;
  LAYER M1 ;
        RECT 14.065 5.795 14.315 6.805 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 4.705 ;
  LAYER M1 ;
        RECT 13.635 7.055 13.885 10.585 ;
  LAYER M1 ;
        RECT 14.495 7.055 14.745 10.585 ;
  LAYER M2 ;
        RECT 13.59 4.06 14.79 4.34 ;
  LAYER M2 ;
        RECT 13.59 9.94 14.79 10.22 ;
  LAYER M2 ;
        RECT 13.16 10.36 14.36 10.64 ;
  LAYER M2 ;
        RECT 13.16 6.16 14.36 6.44 ;
  LAYER M3 ;
        RECT 14.48 4.04 14.76 10.24 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M2 ;
        RECT 8.86 14.14 10.06 14.42 ;
  LAYER M2 ;
        RECT 8.86 7.84 10.06 8.12 ;
  LAYER M2 ;
        RECT 8.86 12.04 10.06 12.32 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M2 ;
        RECT 10.58 0.7 11.78 0.98 ;
  LAYER M2 ;
        RECT 10.58 7 11.78 7.28 ;
  LAYER M2 ;
        RECT 10.58 2.8 11.78 3.08 ;
  LAYER M2 ;
        RECT 11.01 6.58 12.21 6.86 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M2 ;
        RECT 10.58 14.14 11.78 14.42 ;
  LAYER M2 ;
        RECT 10.58 7.84 11.78 8.12 ;
  LAYER M2 ;
        RECT 10.58 12.04 11.78 12.32 ;
  LAYER M2 ;
        RECT 11.01 8.26 12.21 8.54 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M2 ;
        RECT 8.86 0.7 10.06 0.98 ;
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  END 
END TWOBIT_DAC
