* NGSPICE file created from COMPARATOR_0.ext - technology: sky130A
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.subckt NMOS_4T_77406006_X2_Y1_1679747875 a_200_252# a_230_483# a_241_1232# a_147_483#
X0 a_147_483# a_200_252# a_230_483# a_241_1232# sky130_fd_pr__nfet_01v8 ad=6.804e+11p pd=6.66e+06u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X1 a_230_483# a_200_252# a_147_483# a_241_1232# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_147_483# a_200_252# a_230_483# a_241_1232# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_230_483# a_200_252# a_147_483# a_241_1232# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_147_483# a_230_483# 1.31fF
C1 a_200_252# a_230_483# 0.22fF
C2 a_147_483# a_200_252# 0.22fF
C3 a_230_483# a_241_1232# 0.10fF
C4 a_147_483# a_241_1232# 0.32fF
C5 a_200_252# a_241_1232# 1.16fF
.ends

.subckt SCM_PMOS_23436893_X2_Y1_1679747877 a_200_252# a_402_483# w_0_0# VSUBS
X0 w_0_0# a_200_252# a_200_252# w_0_0# sky130_fd_pr__pfet_01v8 ad=1.1508e+12p pd=1.114e+07u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X1 a_402_483# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=0p ps=0u w=840000u l=150000u
X2 a_200_252# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 w_0_0# a_200_252# a_200_252# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 w_0_0# a_200_252# a_402_483# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 a_402_483# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 a_200_252# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 w_0_0# a_200_252# a_402_483# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_402_483# 0.56fF
C1 w_0_0# a_402_483# 1.55fF
C2 a_200_252# w_0_0# 4.37fF
C3 a_402_483# VSUBS -0.14fF
C4 a_200_252# VSUBS 0.04fF
C5 w_0_0# VSUBS 4.49fF
.ends

.subckt NMOS_S_74334133_X2_Y1_1679747876 a_230_483# a_147_483#
X0 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=6.804e+11p pd=6.66e+06u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X1 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_230_483# a_200_252# 0.22fF
C1 a_230_483# a_147_483# 1.46fF
C2 a_200_252# a_147_483# 1.47fF
.ends

.subckt NMOS_S_74334133_X2_Y1_1679747873_1679747874 a_200_252# a_230_483# a_147_483#
X0 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=6.804e+11p pd=6.66e+06u as=4.704e+11p ps=4.48e+06u w=840000u l=150000u
X1 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_230_483# a_200_252# 0.22fF
C1 a_230_483# a_147_483# 1.46fF
C2 a_200_252# a_147_483# 1.47fF
.ends

.subckt PMOS_S_33331942_X2_Y1_1679747874_1679747874 a_200_252# a_230_483# w_0_0# VSUBS
X0 a_230_483# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=4.48e+06u as=6.804e+11p ps=6.66e+06u w=840000u l=150000u
X1 w_0_0# a_200_252# a_230_483# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_230_483# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 w_0_0# a_200_252# a_230_483# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_230_483# 0.22fF
C1 w_0_0# a_230_483# 1.54fF
C2 a_200_252# w_0_0# 1.30fF
C3 a_230_483# VSUBS -0.09fF
C4 a_200_252# VSUBS 0.16fF
C5 w_0_0# VSUBS 3.51fF
.ends

.subckt INV_46031338_PG0_0_0_1679747874 m1_226_560# PMOS_S_33331942_X2_Y1_1679747874_1679747874_0/w_0_0#
+ VSUBS
XNMOS_S_74334133_X2_Y1_1679747873_1679747874_0 m1_226_560# m1_312_1400# VSUBS NMOS_S_74334133_X2_Y1_1679747873_1679747874
XPMOS_S_33331942_X2_Y1_1679747874_1679747874_0 m1_226_560# m1_312_1400# PMOS_S_33331942_X2_Y1_1679747874_1679747874_0/w_0_0#
+ VSUBS PMOS_S_33331942_X2_Y1_1679747874_1679747874
C0 m1_312_1400# PMOS_S_33331942_X2_Y1_1679747874_1679747874_0/w_0_0# 0.02fF
C1 m1_226_560# PMOS_S_33331942_X2_Y1_1679747874_1679747874_0/w_0_0# 0.40fF
C2 m1_226_560# m1_312_1400# 0.27fF
C3 m1_312_1400# VSUBS 1.32fF
C4 m1_226_560# VSUBS 1.86fF
C5 PMOS_S_33331942_X2_Y1_1679747874_1679747874_0/w_0_0# VSUBS 3.59fF
.ends

.subckt COMPARATOR_0
XNMOS_4T_77406006_X2_Y1_1679747875_1 NMOS_4T_77406006_X2_Y1_1679747875_1/a_200_252#
+ m1_602_1400# VSS m1_688_1316# NMOS_4T_77406006_X2_Y1_1679747875
XNMOS_4T_77406006_X2_Y1_1679747875_0 VREF m1_1172_1400# VSS m1_688_1316# NMOS_4T_77406006_X2_Y1_1679747875
XSCM_PMOS_23436893_X2_Y1_1679747877_0 m1_602_1400# m1_1172_1400# VDD VSS SCM_PMOS_23436893_X2_Y1_1679747877
XNMOS_S_74334133_X2_Y1_1679747876_0 m1_688_1316# VSS NMOS_S_74334133_X2_Y1_1679747876
XINV_46031338_PG0_0_0_1679747874_0 m1_1172_1400# VDD VSS INV_46031338_PG0_0_0_1679747874
C0 VREF VIN 0.04fF
C1 OUT VDD 0.16fF
C2 m1_602_1400# VIN 0.00fF
C3 VBIAS m1_1172_1400# 0.00fF
C4 VDD m1_688_1316# 0.26fF
C5 VREF VDD 0.16fF
C6 VBIAS VIN 0.00fF
C7 m1_602_1400# VDD 0.35fF
C8 OUT m1_688_1316# 0.00fF
C9 m1_1172_1400# VIN 0.00fF
C10 OUT m1_602_1400# 0.01fF
C11 VREF m1_688_1316# 0.03fF
C12 VBIAS VDD 0.03fF
C13 m1_602_1400# m1_688_1316# 0.44fF
C14 VREF m1_602_1400# 0.01fF
C15 OUT VBIAS 0.00fF
C16 VDD m1_1172_1400# 0.93fF
C17 OUT m1_1172_1400# 0.01fF
C18 VDD VIN 0.05fF
C19 VBIAS m1_688_1316# 0.00fF
C20 VBIAS m1_602_1400# 0.04fF
C21 m1_1172_1400# m1_688_1316# 0.09fF
C22 VREF m1_1172_1400# 0.04fF
C23 m1_602_1400# m1_1172_1400# 0.39fF
C24 VIN m1_688_1316# 0.01fF
C25 VIN VSS 0.12fF 
C26 VBIAS VSS 0.04fF
C27 OUT VSS 0.12fF 
C28 INV_46031338_PG0_0_0_1679747874_0/m1_312_1400# VSS 1.30fF
C29 m1_1172_1400# VSS 2.08fF
C30 VDD VSS 11.51fF
C31 NMOS_S_74334133_X2_Y1_1679747876_0/a_200_252# VSS 1.47fF $ **FLOATING
C32 m1_688_1316# VSS 1.99fF
C33 VREF VSS 1.14fF
C34 m1_602_1400# VSS 0.07fF
C35 NMOS_4T_77406006_X2_Y1_1679747875_1/a_200_252# VSS 1.16fF
.ends
x1 COMPARATOR_0
V1 VDD VSS 1.8
V2 VIN VSS sine(0 1.8 10000000)
V3 VREF VSS 1
v4 VBIAS VSS 0.9
.tran 10p 10n
.control
run
plot v(VIN) v(VREF) v(VBIAS)
.endc

