MACRO TWO_BIT_DAC
  ORIGIN 0 0 ;
  FOREIGN TWO_BIT_DAC 0 0 ;
  SIZE 31.95 BY 15.71 ;
  PIN D0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.6 2.8 17.8 3.08 ;
      LAYER M2 ;
        RECT 18.32 2.8 19.52 3.08 ;
      LAYER M2 ;
        RECT 17.63 2.8 18.49 3.08 ;
      LAYER M2 ;
        RECT 21.76 2.8 22.96 3.08 ;
      LAYER M2 ;
        RECT 23.48 2.8 24.68 3.08 ;
      LAYER M2 ;
        RECT 22.79 2.8 23.65 3.08 ;
      LAYER M2 ;
        RECT 19.35 2.8 21.93 3.08 ;
    END
  END D0
  PIN X2_INP1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 26.92 7.84 28.12 8.12 ;
      LAYER M3 ;
        RECT 29.96 8.24 30.24 14.44 ;
      LAYER M2 ;
        RECT 27.79 7.84 28.11 8.12 ;
      LAYER M3 ;
        RECT 27.81 7.98 28.09 8.82 ;
      LAYER M2 ;
        RECT 27.95 8.68 30.1 8.96 ;
      LAYER M3 ;
        RECT 29.96 8.635 30.24 9.005 ;
    END
  END X2_INP1
  PIN X2_INP2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 26.92 0.28 28.12 0.56 ;
      LAYER M3 ;
        RECT 29.96 0.68 30.24 6.88 ;
      LAYER M2 ;
        RECT 27.95 0.28 30.1 0.56 ;
      LAYER M3 ;
        RECT 29.96 0.42 30.24 0.84 ;
    END
  END X2_INP2
  PIN X1_INP1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 13.16 7.84 14.36 8.12 ;
      LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
      LAYER M2 ;
        RECT 13.17 7.84 13.49 8.12 ;
      LAYER M3 ;
        RECT 13.19 7.98 13.47 8.82 ;
      LAYER M2 ;
        RECT 11.18 8.68 13.33 8.96 ;
      LAYER M3 ;
        RECT 11.04 8.635 11.32 9.005 ;
    END
  END X1_INP1
  PIN X1_INP2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 13.16 0.28 14.36 0.56 ;
      LAYER M3 ;
        RECT 11.04 0.68 11.32 6.88 ;
      LAYER M2 ;
        RECT 11.18 0.28 13.33 0.56 ;
      LAYER M3 ;
        RECT 11.04 0.42 11.32 0.84 ;
    END
  END X1_INP2
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
      LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
      LAYER M2 ;
        RECT 2.15 12.04 3.01 12.32 ;
    END
  END D1
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 5.88 0.68 6.16 6.88 ;
      LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
      LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
      LAYER M2 ;
        RECT 8.44 7 8.76 7.28 ;
      LAYER M3 ;
        RECT 8.46 7.14 8.74 7.98 ;
      LAYER M2 ;
        RECT 8.44 7.84 8.76 8.12 ;
      LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
      LAYER M3 ;
        RECT 5.88 6.115 6.16 6.485 ;
      LAYER M4 ;
        RECT 6.02 5.9 8.17 6.7 ;
      LAYER M3 ;
        RECT 8.03 6.3 8.31 7.14 ;
      LAYER M2 ;
        RECT 8.01 7 8.33 7.28 ;
      LAYER M3 ;
        RECT 5.88 6.72 6.16 8.4 ;
    END
  END OUT
  OBS 
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M3 ;
        RECT 9.32 14.28 9.6 14.7 ;
  LAYER M2 ;
        RECT 7.31 14.56 9.46 14.84 ;
  LAYER M3 ;
        RECT 26.52 0.68 26.8 6.88 ;
  LAYER M2 ;
        RECT 28.64 7 29.84 7.28 ;
  LAYER M2 ;
        RECT 28.64 7.84 29.84 8.12 ;
  LAYER M2 ;
        RECT 29.08 7 29.4 7.28 ;
  LAYER M3 ;
        RECT 29.1 7.14 29.38 7.98 ;
  LAYER M2 ;
        RECT 29.08 7.84 29.4 8.12 ;
  LAYER M3 ;
        RECT 26.52 8.24 26.8 14.44 ;
  LAYER M3 ;
        RECT 26.52 6.72 26.8 7.14 ;
  LAYER M2 ;
        RECT 26.66 7 28.81 7.28 ;
  LAYER M3 ;
        RECT 26.52 7.14 26.8 8.4 ;
  LAYER M3 ;
        RECT 9.32 9.055 9.6 9.425 ;
  LAYER M2 ;
        RECT 9.46 9.1 26.66 9.38 ;
  LAYER M3 ;
        RECT 26.52 9.055 26.8 9.425 ;
  LAYER M2 ;
        RECT 9.3 9.1 9.62 9.38 ;
  LAYER M3 ;
        RECT 9.32 9.08 9.6 9.4 ;
  LAYER M2 ;
        RECT 26.5 9.1 26.82 9.38 ;
  LAYER M3 ;
        RECT 26.52 9.08 26.8 9.4 ;
  LAYER M2 ;
        RECT 9.3 9.1 9.62 9.38 ;
  LAYER M3 ;
        RECT 9.32 9.08 9.6 9.4 ;
  LAYER M2 ;
        RECT 26.5 9.1 26.82 9.38 ;
  LAYER M3 ;
        RECT 26.52 9.08 26.8 9.4 ;
  LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M3 ;
        RECT 9.32 6.115 9.6 6.485 ;
  LAYER M2 ;
        RECT 7.31 6.16 9.46 6.44 ;
  LAYER M1 ;
        RECT 7.185 6.3 7.435 7.14 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 14.48 0.68 14.76 6.88 ;
  LAYER M2 ;
        RECT 11.44 7 12.64 7.28 ;
  LAYER M2 ;
        RECT 11.44 7.84 12.64 8.12 ;
  LAYER M2 ;
        RECT 11.88 7 12.2 7.28 ;
  LAYER M3 ;
        RECT 11.9 7.14 12.18 7.98 ;
  LAYER M2 ;
        RECT 11.88 7.84 12.2 8.12 ;
  LAYER M3 ;
        RECT 14.48 8.24 14.76 14.44 ;
  LAYER M3 ;
        RECT 14.48 6.72 14.76 7.14 ;
  LAYER M2 ;
        RECT 12.47 7 14.62 7.28 ;
  LAYER M3 ;
        RECT 14.48 7.14 14.76 8.4 ;
  LAYER M2 ;
        RECT 9.46 6.16 11.61 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.3 11.75 7.14 ;
  LAYER M2 ;
        RECT 11.45 7 11.77 7.28 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M2 ;
        RECT 11.45 7 11.77 7.28 ;
  LAYER M3 ;
        RECT 11.47 6.98 11.75 7.3 ;
  LAYER M2 ;
        RECT 11.45 6.16 11.77 6.44 ;
  LAYER M3 ;
        RECT 11.47 6.14 11.75 6.46 ;
  LAYER M2 ;
        RECT 11.45 7 11.77 7.28 ;
  LAYER M3 ;
        RECT 11.47 6.98 11.75 7.3 ;
  LAYER M2 ;
        RECT 21.76 7.84 22.96 8.12 ;
  LAYER M2 ;
        RECT 24.34 7.84 25.54 8.12 ;
  LAYER M2 ;
        RECT 28.64 2.8 29.84 3.08 ;
  LAYER M2 ;
        RECT 28.64 12.04 29.84 12.32 ;
  LAYER M2 ;
        RECT 28.65 2.8 28.97 3.08 ;
  LAYER M1 ;
        RECT 28.685 2.94 28.935 12.18 ;
  LAYER M2 ;
        RECT 28.65 12.04 28.97 12.32 ;
  LAYER M2 ;
        RECT 22.79 7.84 24.51 8.12 ;
  LAYER M2 ;
        RECT 25.37 7.84 26.23 8.12 ;
  LAYER M1 ;
        RECT 26.105 7.56 26.355 7.98 ;
  LAYER M2 ;
        RECT 26.23 7.42 28.81 7.7 ;
  LAYER M1 ;
        RECT 28.685 7.475 28.935 7.645 ;
  LAYER M1 ;
        RECT 26.105 7.475 26.355 7.645 ;
  LAYER M2 ;
        RECT 26.06 7.42 26.4 7.7 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 8.065 ;
  LAYER M2 ;
        RECT 26.06 7.84 26.4 8.12 ;
  LAYER M1 ;
        RECT 28.685 7.475 28.935 7.645 ;
  LAYER M2 ;
        RECT 28.64 7.42 28.98 7.7 ;
  LAYER M1 ;
        RECT 26.105 7.475 26.355 7.645 ;
  LAYER M2 ;
        RECT 26.06 7.42 26.4 7.7 ;
  LAYER M1 ;
        RECT 26.105 7.895 26.355 8.065 ;
  LAYER M2 ;
        RECT 26.06 7.84 26.4 8.12 ;
  LAYER M1 ;
        RECT 28.685 7.475 28.935 7.645 ;
  LAYER M2 ;
        RECT 28.64 7.42 28.98 7.7 ;
  LAYER M2 ;
        RECT 21.76 7 22.96 7.28 ;
  LAYER M2 ;
        RECT 23.48 7 24.68 7.28 ;
  LAYER M2 ;
        RECT 21.76 12.04 22.96 12.32 ;
  LAYER M2 ;
        RECT 24.34 12.04 25.54 12.32 ;
  LAYER M2 ;
        RECT 26.92 12.04 28.12 12.32 ;
  LAYER M2 ;
        RECT 26.92 4.48 28.12 4.76 ;
  LAYER M2 ;
        RECT 22.79 7 23.65 7.28 ;
  LAYER M2 ;
        RECT 22.63 7 22.95 7.28 ;
  LAYER M1 ;
        RECT 22.665 7.14 22.915 12.18 ;
  LAYER M2 ;
        RECT 22.63 12.04 22.95 12.32 ;
  LAYER M2 ;
        RECT 22.79 12.04 24.51 12.32 ;
  LAYER M2 ;
        RECT 25.37 12.04 27.09 12.32 ;
  LAYER M2 ;
        RECT 24.35 7 24.67 7.28 ;
  LAYER M3 ;
        RECT 24.37 4.62 24.65 7.14 ;
  LAYER M2 ;
        RECT 24.51 4.48 27.09 4.76 ;
  LAYER M1 ;
        RECT 22.665 7.055 22.915 7.225 ;
  LAYER M2 ;
        RECT 22.62 7 22.96 7.28 ;
  LAYER M1 ;
        RECT 22.665 12.095 22.915 12.265 ;
  LAYER M2 ;
        RECT 22.62 12.04 22.96 12.32 ;
  LAYER M1 ;
        RECT 22.665 7.055 22.915 7.225 ;
  LAYER M2 ;
        RECT 22.62 7 22.96 7.28 ;
  LAYER M1 ;
        RECT 22.665 12.095 22.915 12.265 ;
  LAYER M2 ;
        RECT 22.62 12.04 22.96 12.32 ;
  LAYER M1 ;
        RECT 22.665 7.055 22.915 7.225 ;
  LAYER M2 ;
        RECT 22.62 7 22.96 7.28 ;
  LAYER M1 ;
        RECT 22.665 12.095 22.915 12.265 ;
  LAYER M2 ;
        RECT 22.62 12.04 22.96 12.32 ;
  LAYER M1 ;
        RECT 22.665 7.055 22.915 7.225 ;
  LAYER M2 ;
        RECT 22.62 7 22.96 7.28 ;
  LAYER M1 ;
        RECT 22.665 12.095 22.915 12.265 ;
  LAYER M2 ;
        RECT 22.62 12.04 22.96 12.32 ;
  LAYER M1 ;
        RECT 22.665 7.055 22.915 7.225 ;
  LAYER M2 ;
        RECT 22.62 7 22.96 7.28 ;
  LAYER M1 ;
        RECT 22.665 12.095 22.915 12.265 ;
  LAYER M2 ;
        RECT 22.62 12.04 22.96 12.32 ;
  LAYER M1 ;
        RECT 22.665 7.055 22.915 7.225 ;
  LAYER M2 ;
        RECT 22.62 7 22.96 7.28 ;
  LAYER M1 ;
        RECT 22.665 12.095 22.915 12.265 ;
  LAYER M2 ;
        RECT 22.62 12.04 22.96 12.32 ;
  LAYER M1 ;
        RECT 22.665 7.055 22.915 7.225 ;
  LAYER M2 ;
        RECT 22.62 7 22.96 7.28 ;
  LAYER M1 ;
        RECT 22.665 12.095 22.915 12.265 ;
  LAYER M2 ;
        RECT 22.62 12.04 22.96 12.32 ;
  LAYER M2 ;
        RECT 24.35 4.48 24.67 4.76 ;
  LAYER M3 ;
        RECT 24.37 4.46 24.65 4.78 ;
  LAYER M2 ;
        RECT 24.35 7 24.67 7.28 ;
  LAYER M3 ;
        RECT 24.37 6.98 24.65 7.3 ;
  LAYER M1 ;
        RECT 22.665 7.055 22.915 7.225 ;
  LAYER M2 ;
        RECT 22.62 7 22.96 7.28 ;
  LAYER M1 ;
        RECT 22.665 12.095 22.915 12.265 ;
  LAYER M2 ;
        RECT 22.62 12.04 22.96 12.32 ;
  LAYER M2 ;
        RECT 24.35 4.48 24.67 4.76 ;
  LAYER M3 ;
        RECT 24.37 4.46 24.65 4.78 ;
  LAYER M2 ;
        RECT 24.35 7 24.67 7.28 ;
  LAYER M3 ;
        RECT 24.37 6.98 24.65 7.3 ;
  LAYER M1 ;
        RECT 29.545 3.695 29.795 7.225 ;
  LAYER M1 ;
        RECT 29.545 2.435 29.795 3.445 ;
  LAYER M1 ;
        RECT 29.545 0.335 29.795 1.345 ;
  LAYER M1 ;
        RECT 29.115 3.695 29.365 7.225 ;
  LAYER M1 ;
        RECT 29.975 3.695 30.225 7.225 ;
  LAYER M2 ;
        RECT 29.07 0.7 30.27 0.98 ;
  LAYER M2 ;
        RECT 29.07 6.58 30.27 6.86 ;
  LAYER M2 ;
        RECT 28.64 7 29.84 7.28 ;
  LAYER M2 ;
        RECT 28.64 2.8 29.84 3.08 ;
  LAYER M3 ;
        RECT 29.96 0.68 30.24 6.88 ;
  LAYER M1 ;
        RECT 29.545 7.895 29.795 11.425 ;
  LAYER M1 ;
        RECT 29.545 11.675 29.795 12.685 ;
  LAYER M1 ;
        RECT 29.545 13.775 29.795 14.785 ;
  LAYER M1 ;
        RECT 29.115 7.895 29.365 11.425 ;
  LAYER M1 ;
        RECT 29.975 7.895 30.225 11.425 ;
  LAYER M2 ;
        RECT 29.07 14.14 30.27 14.42 ;
  LAYER M2 ;
        RECT 29.07 8.26 30.27 8.54 ;
  LAYER M2 ;
        RECT 28.64 7.84 29.84 8.12 ;
  LAYER M2 ;
        RECT 28.64 12.04 29.84 12.32 ;
  LAYER M3 ;
        RECT 29.96 8.24 30.24 14.44 ;
  LAYER M1 ;
        RECT 21.805 3.695 22.055 7.225 ;
  LAYER M1 ;
        RECT 21.805 2.435 22.055 3.445 ;
  LAYER M1 ;
        RECT 21.805 0.335 22.055 1.345 ;
  LAYER M1 ;
        RECT 22.235 3.695 22.485 7.225 ;
  LAYER M1 ;
        RECT 21.375 3.695 21.625 7.225 ;
  LAYER M2 ;
        RECT 21.33 0.7 22.53 0.98 ;
  LAYER M2 ;
        RECT 21.33 6.58 22.53 6.86 ;
  LAYER M2 ;
        RECT 21.76 7 22.96 7.28 ;
  LAYER M2 ;
        RECT 21.76 2.8 22.96 3.08 ;
  LAYER M3 ;
        RECT 21.36 0.68 21.64 6.88 ;
  LAYER M1 ;
        RECT 24.385 7.895 24.635 11.425 ;
  LAYER M1 ;
        RECT 24.385 11.675 24.635 12.685 ;
  LAYER M1 ;
        RECT 24.385 13.775 24.635 14.785 ;
  LAYER M1 ;
        RECT 24.815 7.895 25.065 11.425 ;
  LAYER M1 ;
        RECT 23.955 7.895 24.205 11.425 ;
  LAYER M2 ;
        RECT 23.91 14.14 25.11 14.42 ;
  LAYER M2 ;
        RECT 23.91 8.26 25.11 8.54 ;
  LAYER M2 ;
        RECT 24.34 7.84 25.54 8.12 ;
  LAYER M2 ;
        RECT 24.34 12.04 25.54 12.32 ;
  LAYER M3 ;
        RECT 23.94 8.24 24.22 14.44 ;
  LAYER M1 ;
        RECT 26.965 7.895 27.215 11.425 ;
  LAYER M1 ;
        RECT 26.965 11.675 27.215 12.685 ;
  LAYER M1 ;
        RECT 26.965 13.775 27.215 14.785 ;
  LAYER M1 ;
        RECT 27.395 7.895 27.645 11.425 ;
  LAYER M1 ;
        RECT 26.535 7.895 26.785 11.425 ;
  LAYER M2 ;
        RECT 26.49 14.14 27.69 14.42 ;
  LAYER M2 ;
        RECT 26.49 8.26 27.69 8.54 ;
  LAYER M2 ;
        RECT 26.92 7.84 28.12 8.12 ;
  LAYER M2 ;
        RECT 26.92 12.04 28.12 12.32 ;
  LAYER M3 ;
        RECT 26.52 8.24 26.8 14.44 ;
  LAYER M1 ;
        RECT 24.385 3.695 24.635 7.225 ;
  LAYER M1 ;
        RECT 24.385 2.435 24.635 3.445 ;
  LAYER M1 ;
        RECT 24.385 0.335 24.635 1.345 ;
  LAYER M1 ;
        RECT 23.955 3.695 24.205 7.225 ;
  LAYER M1 ;
        RECT 24.815 3.695 25.065 7.225 ;
  LAYER M2 ;
        RECT 23.91 0.7 25.11 0.98 ;
  LAYER M2 ;
        RECT 23.91 6.58 25.11 6.86 ;
  LAYER M2 ;
        RECT 23.48 7 24.68 7.28 ;
  LAYER M2 ;
        RECT 23.48 2.8 24.68 3.08 ;
  LAYER M3 ;
        RECT 24.8 0.68 25.08 6.88 ;
  LAYER M1 ;
        RECT 21.805 7.895 22.055 11.425 ;
  LAYER M1 ;
        RECT 21.805 11.675 22.055 12.685 ;
  LAYER M1 ;
        RECT 21.805 13.775 22.055 14.785 ;
  LAYER M1 ;
        RECT 22.235 7.895 22.485 11.425 ;
  LAYER M1 ;
        RECT 21.375 7.895 21.625 11.425 ;
  LAYER M2 ;
        RECT 21.33 14.14 22.53 14.42 ;
  LAYER M2 ;
        RECT 21.33 8.26 22.53 8.54 ;
  LAYER M2 ;
        RECT 21.76 7.84 22.96 8.12 ;
  LAYER M2 ;
        RECT 21.76 12.04 22.96 12.32 ;
  LAYER M3 ;
        RECT 21.36 8.24 21.64 14.44 ;
  LAYER M1 ;
        RECT 26.965 0.335 27.215 3.865 ;
  LAYER M1 ;
        RECT 26.965 4.115 27.215 5.125 ;
  LAYER M1 ;
        RECT 26.965 6.215 27.215 7.225 ;
  LAYER M1 ;
        RECT 27.395 0.335 27.645 3.865 ;
  LAYER M1 ;
        RECT 26.535 0.335 26.785 3.865 ;
  LAYER M2 ;
        RECT 26.49 6.58 27.69 6.86 ;
  LAYER M2 ;
        RECT 26.49 0.7 27.69 0.98 ;
  LAYER M2 ;
        RECT 26.92 0.28 28.12 0.56 ;
  LAYER M2 ;
        RECT 26.92 4.48 28.12 4.76 ;
  LAYER M3 ;
        RECT 26.52 0.68 26.8 6.88 ;
  LAYER M2 ;
        RECT 11.44 2.8 12.64 3.08 ;
  LAYER M2 ;
        RECT 11.44 12.04 12.64 12.32 ;
  LAYER M2 ;
        RECT 12.31 2.8 12.63 3.08 ;
  LAYER M1 ;
        RECT 12.345 2.94 12.595 12.18 ;
  LAYER M2 ;
        RECT 12.31 12.04 12.63 12.32 ;
  LAYER M2 ;
        RECT 15.74 7.84 16.94 8.12 ;
  LAYER M2 ;
        RECT 18.32 7.84 19.52 8.12 ;
  LAYER M1 ;
        RECT 12.345 7.475 12.595 7.645 ;
  LAYER M2 ;
        RECT 12.47 7.42 15.05 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.56 15.175 7.98 ;
  LAYER M2 ;
        RECT 15.05 7.84 15.91 8.12 ;
  LAYER M2 ;
        RECT 16.77 7.84 18.49 8.12 ;
  LAYER M1 ;
        RECT 12.345 7.475 12.595 7.645 ;
  LAYER M2 ;
        RECT 12.3 7.42 12.64 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.475 15.175 7.645 ;
  LAYER M2 ;
        RECT 14.88 7.42 15.22 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 8.065 ;
  LAYER M2 ;
        RECT 14.88 7.84 15.22 8.12 ;
  LAYER M1 ;
        RECT 12.345 7.475 12.595 7.645 ;
  LAYER M2 ;
        RECT 12.3 7.42 12.64 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.475 15.175 7.645 ;
  LAYER M2 ;
        RECT 14.88 7.42 15.22 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 8.065 ;
  LAYER M2 ;
        RECT 14.88 7.84 15.22 8.12 ;
  LAYER M1 ;
        RECT 12.345 7.475 12.595 7.645 ;
  LAYER M2 ;
        RECT 12.3 7.42 12.64 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.475 15.175 7.645 ;
  LAYER M2 ;
        RECT 14.88 7.42 15.22 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 8.065 ;
  LAYER M2 ;
        RECT 14.88 7.84 15.22 8.12 ;
  LAYER M1 ;
        RECT 12.345 7.475 12.595 7.645 ;
  LAYER M2 ;
        RECT 12.3 7.42 12.64 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.475 15.175 7.645 ;
  LAYER M2 ;
        RECT 14.88 7.42 15.22 7.7 ;
  LAYER M1 ;
        RECT 14.925 7.895 15.175 8.065 ;
  LAYER M2 ;
        RECT 14.88 7.84 15.22 8.12 ;
  LAYER M2 ;
        RECT 13.16 4.48 14.36 4.76 ;
  LAYER M2 ;
        RECT 16.6 7 17.8 7.28 ;
  LAYER M2 ;
        RECT 18.32 7 19.52 7.28 ;
  LAYER M2 ;
        RECT 18.32 12.04 19.52 12.32 ;
  LAYER M2 ;
        RECT 15.74 12.04 16.94 12.32 ;
  LAYER M2 ;
        RECT 13.16 12.04 14.36 12.32 ;
  LAYER M2 ;
        RECT 14.19 4.48 16.77 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.62 16.91 7.14 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M2 ;
        RECT 17.63 7 18.49 7.28 ;
  LAYER M2 ;
        RECT 18.33 7 18.65 7.28 ;
  LAYER M1 ;
        RECT 18.365 7.14 18.615 12.18 ;
  LAYER M2 ;
        RECT 18.33 12.04 18.65 12.32 ;
  LAYER M2 ;
        RECT 16.77 12.04 18.49 12.32 ;
  LAYER M2 ;
        RECT 14.19 12.04 15.91 12.32 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M1 ;
        RECT 18.365 7.055 18.615 7.225 ;
  LAYER M2 ;
        RECT 18.32 7 18.66 7.28 ;
  LAYER M1 ;
        RECT 18.365 12.095 18.615 12.265 ;
  LAYER M2 ;
        RECT 18.32 12.04 18.66 12.32 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M1 ;
        RECT 18.365 7.055 18.615 7.225 ;
  LAYER M2 ;
        RECT 18.32 7 18.66 7.28 ;
  LAYER M1 ;
        RECT 18.365 12.095 18.615 12.265 ;
  LAYER M2 ;
        RECT 18.32 12.04 18.66 12.32 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M1 ;
        RECT 18.365 7.055 18.615 7.225 ;
  LAYER M2 ;
        RECT 18.32 7 18.66 7.28 ;
  LAYER M1 ;
        RECT 18.365 12.095 18.615 12.265 ;
  LAYER M2 ;
        RECT 18.32 12.04 18.66 12.32 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M1 ;
        RECT 18.365 7.055 18.615 7.225 ;
  LAYER M2 ;
        RECT 18.32 7 18.66 7.28 ;
  LAYER M1 ;
        RECT 18.365 12.095 18.615 12.265 ;
  LAYER M2 ;
        RECT 18.32 12.04 18.66 12.32 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M1 ;
        RECT 18.365 7.055 18.615 7.225 ;
  LAYER M2 ;
        RECT 18.32 7 18.66 7.28 ;
  LAYER M1 ;
        RECT 18.365 12.095 18.615 12.265 ;
  LAYER M2 ;
        RECT 18.32 12.04 18.66 12.32 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M1 ;
        RECT 18.365 7.055 18.615 7.225 ;
  LAYER M2 ;
        RECT 18.32 7 18.66 7.28 ;
  LAYER M1 ;
        RECT 18.365 12.095 18.615 12.265 ;
  LAYER M2 ;
        RECT 18.32 12.04 18.66 12.32 ;
  LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
  LAYER M3 ;
        RECT 16.63 4.46 16.91 4.78 ;
  LAYER M2 ;
        RECT 16.61 7 16.93 7.28 ;
  LAYER M3 ;
        RECT 16.63 6.98 16.91 7.3 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M2 ;
        RECT 11.01 0.7 12.21 0.98 ;
  LAYER M2 ;
        RECT 11.01 6.58 12.21 6.86 ;
  LAYER M2 ;
        RECT 11.44 7 12.64 7.28 ;
  LAYER M2 ;
        RECT 11.44 2.8 12.64 3.08 ;
  LAYER M3 ;
        RECT 11.04 0.68 11.32 6.88 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 11.425 ;
  LAYER M1 ;
        RECT 11.485 11.675 11.735 12.685 ;
  LAYER M1 ;
        RECT 11.485 13.775 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.915 7.895 12.165 11.425 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M2 ;
        RECT 11.01 14.14 12.21 14.42 ;
  LAYER M2 ;
        RECT 11.01 8.26 12.21 8.54 ;
  LAYER M2 ;
        RECT 11.44 7.84 12.64 8.12 ;
  LAYER M2 ;
        RECT 11.44 12.04 12.64 12.32 ;
  LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
  LAYER M1 ;
        RECT 19.225 3.695 19.475 7.225 ;
  LAYER M1 ;
        RECT 19.225 2.435 19.475 3.445 ;
  LAYER M1 ;
        RECT 19.225 0.335 19.475 1.345 ;
  LAYER M1 ;
        RECT 18.795 3.695 19.045 7.225 ;
  LAYER M1 ;
        RECT 19.655 3.695 19.905 7.225 ;
  LAYER M2 ;
        RECT 18.75 0.7 19.95 0.98 ;
  LAYER M2 ;
        RECT 18.75 6.58 19.95 6.86 ;
  LAYER M2 ;
        RECT 18.32 7 19.52 7.28 ;
  LAYER M2 ;
        RECT 18.32 2.8 19.52 3.08 ;
  LAYER M3 ;
        RECT 19.64 0.68 19.92 6.88 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 12.685 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 14.785 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M2 ;
        RECT 16.17 14.14 17.37 14.42 ;
  LAYER M2 ;
        RECT 16.17 8.26 17.37 8.54 ;
  LAYER M2 ;
        RECT 15.74 7.84 16.94 8.12 ;
  LAYER M2 ;
        RECT 15.74 12.04 16.94 12.32 ;
  LAYER M3 ;
        RECT 17.06 8.24 17.34 14.44 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M2 ;
        RECT 13.59 14.14 14.79 14.42 ;
  LAYER M2 ;
        RECT 13.59 8.26 14.79 8.54 ;
  LAYER M2 ;
        RECT 13.16 7.84 14.36 8.12 ;
  LAYER M2 ;
        RECT 13.16 12.04 14.36 12.32 ;
  LAYER M3 ;
        RECT 14.48 8.24 14.76 14.44 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M2 ;
        RECT 16.17 0.7 17.37 0.98 ;
  LAYER M2 ;
        RECT 16.17 6.58 17.37 6.86 ;
  LAYER M2 ;
        RECT 16.6 7 17.8 7.28 ;
  LAYER M2 ;
        RECT 16.6 2.8 17.8 3.08 ;
  LAYER M3 ;
        RECT 16.2 0.68 16.48 6.88 ;
  LAYER M1 ;
        RECT 19.225 7.895 19.475 11.425 ;
  LAYER M1 ;
        RECT 19.225 11.675 19.475 12.685 ;
  LAYER M1 ;
        RECT 19.225 13.775 19.475 14.785 ;
  LAYER M1 ;
        RECT 18.795 7.895 19.045 11.425 ;
  LAYER M1 ;
        RECT 19.655 7.895 19.905 11.425 ;
  LAYER M2 ;
        RECT 18.75 14.14 19.95 14.42 ;
  LAYER M2 ;
        RECT 18.75 8.26 19.95 8.54 ;
  LAYER M2 ;
        RECT 18.32 7.84 19.52 8.12 ;
  LAYER M2 ;
        RECT 18.32 12.04 19.52 12.32 ;
  LAYER M3 ;
        RECT 19.64 8.24 19.92 14.44 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 3.865 ;
  LAYER M1 ;
        RECT 14.065 4.115 14.315 5.125 ;
  LAYER M1 ;
        RECT 14.065 6.215 14.315 7.225 ;
  LAYER M1 ;
        RECT 13.635 0.335 13.885 3.865 ;
  LAYER M1 ;
        RECT 14.495 0.335 14.745 3.865 ;
  LAYER M2 ;
        RECT 13.59 6.58 14.79 6.86 ;
  LAYER M2 ;
        RECT 13.59 0.7 14.79 0.98 ;
  LAYER M2 ;
        RECT 13.16 0.28 14.36 0.56 ;
  LAYER M2 ;
        RECT 13.16 4.48 14.36 4.76 ;
  LAYER M3 ;
        RECT 14.48 0.68 14.76 6.88 ;
  LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M2 ;
        RECT 8.01 2.8 8.33 3.08 ;
  LAYER M1 ;
        RECT 8.045 2.94 8.295 12.18 ;
  LAYER M2 ;
        RECT 8.01 12.04 8.33 12.32 ;
  LAYER M2 ;
        RECT 2.15 7 3.87 7.28 ;
  LAYER M2 ;
        RECT 4.73 7 5.59 7.28 ;
  LAYER M1 ;
        RECT 5.465 7.14 5.715 7.56 ;
  LAYER M2 ;
        RECT 5.59 7.42 8.17 7.7 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M1 ;
        RECT 5.465 7.055 5.715 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 5.76 7.28 ;
  LAYER M1 ;
        RECT 5.465 7.475 5.715 7.645 ;
  LAYER M2 ;
        RECT 5.42 7.42 5.76 7.7 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M2 ;
        RECT 8 7.42 8.34 7.7 ;
  LAYER M1 ;
        RECT 5.465 7.055 5.715 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 5.76 7.28 ;
  LAYER M1 ;
        RECT 5.465 7.475 5.715 7.645 ;
  LAYER M2 ;
        RECT 5.42 7.42 5.76 7.7 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M2 ;
        RECT 8 7.42 8.34 7.7 ;
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
  LAYER M2 ;
        RECT 2.15 2.8 3.87 3.08 ;
  LAYER M2 ;
        RECT 4.73 2.8 6.45 3.08 ;
  LAYER M2 ;
        RECT 1.99 2.8 2.31 3.08 ;
  LAYER M1 ;
        RECT 2.025 2.94 2.275 7.98 ;
  LAYER M2 ;
        RECT 1.99 7.84 2.31 8.12 ;
  LAYER M2 ;
        RECT 2.15 7.84 3.01 8.12 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.98 4.01 10.5 ;
  LAYER M2 ;
        RECT 3.87 10.36 6.45 10.64 ;
  LAYER M1 ;
        RECT 2.025 2.855 2.275 3.025 ;
  LAYER M2 ;
        RECT 1.98 2.8 2.32 3.08 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 2.855 2.275 3.025 ;
  LAYER M2 ;
        RECT 1.98 2.8 2.32 3.08 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 2.855 2.275 3.025 ;
  LAYER M2 ;
        RECT 1.98 2.8 2.32 3.08 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 2.855 2.275 3.025 ;
  LAYER M2 ;
        RECT 1.98 2.8 2.32 3.08 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 2.855 2.275 3.025 ;
  LAYER M2 ;
        RECT 1.98 2.8 2.32 3.08 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M2 ;
        RECT 3.71 10.36 4.03 10.64 ;
  LAYER M3 ;
        RECT 3.73 10.34 4.01 10.66 ;
  LAYER M1 ;
        RECT 2.025 2.855 2.275 3.025 ;
  LAYER M2 ;
        RECT 1.98 2.8 2.32 3.08 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M2 ;
        RECT 3.71 10.36 4.03 10.64 ;
  LAYER M3 ;
        RECT 3.73 10.34 4.01 10.66 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M2 ;
        RECT 8.43 14.14 9.63 14.42 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M3 ;
        RECT 0.72 8.24 1 14.44 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M2 ;
        RECT 5.85 6.58 7.05 6.86 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 6.88 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M3 ;
        RECT 0.72 0.68 1 6.88 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
  END 
END TWO_BIT_DAC
