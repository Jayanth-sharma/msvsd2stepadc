* SPICE3 file created from INVERTER_0.ext - technology: sky130A
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

x1 A B VDD VSS inverter



.subckt inverter A B VDD VSS
X0 B A VSS VSS sky130_fd_pr__nfet_01v8 ad=2.94e+12p pd=2.38e+07u as=3.465e+12p ps=2.85e+07u w=2.1e+06u l=150000u
X1 VSS A B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X2 B A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X3 VSS A B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X4 VSS A B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X5 B A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X6 B A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X7 VSS A B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X8 VSS A B VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X9 B A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X10 B A INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+12p pd=2.38e+07u as=3.465e+12p ps=2.85e+07u w=2.1e+06u l=150000u
X11 INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# A B INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X12 INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# A B INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X13 B A INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X14 B A INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X15 INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# A B INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X16 INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# A B INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X17 B A INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X18 B A INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X19 INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# A B INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
C0 B A 1.20fF
C1 INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# A 2.60fF
C2 INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# B 4.03fF
C3 B VSS 3.35fF 
C4 A VSS 2.98fF 
C5 INV_986780_0_0_1677685626_0/PMOS_S_86637345_X5_Y1_1677685627_1677685626_0/w_0_0# VSS 5.63fF 

.ends
Vgnd VSS 0 0 
VDD VDD VSS 1.8
Vin A  VSS 0
* create pulse 
* Vin A VSS pulse(0 1.8 1p 10p 10p 1n 2n)

* create PWL 
* Vin A VSS pwl(0 1.8v 5n 1.8v 5.1n 0 10n 0)
* .tran 10p 10n


.dc Vin 0 1.8 0.01


.control
  run 
  plot A B
.endc 

.end

