magic
tech sky130A
magscale 1 2
timestamp 1679679491
<< locali >>
rect 577 1831 585 1865
rect 619 1831 627 1865
rect 405 1747 413 1781
rect 447 1747 455 1781
rect 577 17 627 1831
rect 577 -17 585 17
rect 619 -17 627 17
rect 1437 1747 1445 1781
rect 1479 1747 1487 1781
rect 1437 17 1487 1747
rect 1437 -17 1445 17
rect 1479 -17 1487 17
<< viali >>
rect 585 1831 619 1865
rect 413 1747 447 1781
rect 585 -17 619 17
rect 1445 1747 1479 1781
rect 1445 -17 1479 17
<< metal1 >>
rect 568 1874 720 1876
rect 568 1865 662 1874
rect 568 1831 585 1865
rect 619 1831 662 1865
rect 568 1822 662 1831
rect 714 1822 720 1874
rect 568 1820 720 1822
rect 140 1790 290 1792
rect 140 1738 146 1790
rect 198 1738 232 1790
rect 284 1738 290 1790
rect 140 1736 290 1738
rect 396 1790 1150 1792
rect 396 1781 1092 1790
rect 396 1747 413 1781
rect 447 1747 1092 1781
rect 396 1738 1092 1747
rect 1144 1738 1150 1790
rect 396 1736 1150 1738
rect 1344 1790 1496 1792
rect 1344 1738 1350 1790
rect 1402 1781 1496 1790
rect 1402 1747 1445 1781
rect 1479 1747 1496 1781
rect 1402 1738 1496 1747
rect 1344 1736 1496 1738
rect 1086 1622 1150 1624
rect 1086 1570 1092 1622
rect 1144 1570 1150 1622
rect 1086 1568 1150 1570
rect 312 1538 892 1540
rect 312 1486 318 1538
rect 370 1486 834 1538
rect 886 1486 892 1538
rect 312 1484 892 1486
rect 54 1286 204 1288
rect 54 1234 60 1286
rect 112 1234 146 1286
rect 198 1234 204 1286
rect 54 1232 204 1234
rect 570 1286 720 1288
rect 570 1234 576 1286
rect 628 1234 662 1286
rect 714 1234 720 1286
rect 570 1232 720 1234
rect 1258 1286 1408 1288
rect 1258 1234 1264 1286
rect 1316 1234 1350 1286
rect 1402 1234 1408 1286
rect 1258 1232 1408 1234
rect 568 26 636 28
rect 568 -26 576 26
rect 628 -26 636 26
rect 568 -28 636 -26
rect 1258 26 1496 28
rect 1258 -26 1264 26
rect 1316 17 1496 26
rect 1316 -17 1445 17
rect 1479 -17 1496 17
rect 1316 -26 1496 -17
rect 1258 -28 1496 -26
<< via1 >>
rect 662 1822 714 1874
rect 146 1738 198 1790
rect 232 1738 284 1790
rect 1092 1738 1144 1790
rect 1350 1738 1402 1790
rect 1092 1570 1144 1622
rect 318 1486 370 1538
rect 834 1486 886 1538
rect 60 1234 112 1286
rect 146 1234 198 1286
rect 576 1234 628 1286
rect 662 1234 714 1286
rect 1264 1234 1316 1286
rect 1350 1234 1402 1286
rect 576 17 628 26
rect 576 -17 585 17
rect 585 -17 619 17
rect 619 -17 628 17
rect 576 -26 628 -17
rect 1264 -26 1316 26
<< metal2 >>
rect 660 1874 716 1880
rect 660 1822 662 1874
rect 714 1822 716 1874
rect 660 1816 716 1822
rect 58 1792 114 1801
rect 58 1286 114 1736
rect 144 1790 200 1796
rect 144 1738 146 1790
rect 198 1738 200 1790
rect 144 1732 200 1738
rect 230 1790 286 1796
rect 230 1738 232 1790
rect 284 1738 286 1790
rect 58 1234 60 1286
rect 112 1234 114 1286
rect 58 1228 114 1234
rect 144 1286 200 1292
rect 144 1234 146 1286
rect 198 1234 200 1286
rect 144 1228 200 1234
rect 230 28 286 1738
rect 574 1792 630 1801
rect 316 1538 372 1544
rect 316 1486 318 1538
rect 370 1486 372 1538
rect 316 1480 372 1486
rect 574 1286 630 1736
rect 1090 1790 1146 1796
rect 1090 1738 1092 1790
rect 1144 1738 1146 1790
rect 1090 1622 1146 1738
rect 1090 1570 1092 1622
rect 1144 1570 1146 1622
rect 1090 1564 1146 1570
rect 1262 1792 1318 1801
rect 832 1538 888 1544
rect 832 1486 834 1538
rect 886 1486 888 1538
rect 832 1480 888 1486
rect 574 1234 576 1286
rect 628 1234 630 1286
rect 574 1228 630 1234
rect 660 1286 716 1292
rect 660 1234 662 1286
rect 714 1234 716 1286
rect 660 1228 716 1234
rect 1262 1286 1318 1736
rect 1348 1790 1404 1796
rect 1348 1738 1350 1790
rect 1402 1738 1404 1790
rect 1348 1732 1404 1738
rect 1262 1234 1264 1286
rect 1316 1234 1318 1286
rect 1262 1228 1318 1234
rect 1348 1286 1404 1292
rect 1348 1234 1350 1286
rect 1402 1234 1404 1286
rect 1348 1228 1404 1234
rect 230 -37 286 -28
rect 574 28 630 48
rect 574 -37 630 -28
rect 1262 28 1318 48
rect 1262 -37 1318 -28
<< via2 >>
rect 58 1736 114 1792
rect 574 1736 630 1792
rect 1262 1736 1318 1792
rect 230 -28 286 28
rect 574 26 630 28
rect 574 -26 576 26
rect 576 -26 628 26
rect 628 -26 630 26
rect 574 -28 630 -26
rect 1262 26 1318 28
rect 1262 -26 1264 26
rect 1264 -26 1316 26
rect 1316 -26 1318 26
rect 1262 -28 1318 -26
<< metal3 >>
rect -80 1796 2448 1844
rect -80 1792 2336 1796
rect -80 1736 58 1792
rect 114 1736 574 1792
rect 630 1736 1262 1792
rect 1318 1736 2336 1792
rect -80 1732 2336 1736
rect 2400 1732 2448 1796
rect -80 1684 2448 1732
rect -80 32 2448 80
rect -80 -32 -32 32
rect 32 28 2448 32
rect 32 -28 230 28
rect 286 -28 574 28
rect 630 -28 1262 28
rect 1318 -28 2448 28
rect 32 -32 2448 -28
rect -80 -80 2448 -32
<< via3 >>
rect 2336 1732 2400 1796
rect -32 -32 32 32
<< metal4 >>
rect -118 32 118 1882
rect -118 -32 -32 32
rect 32 -32 118 32
rect -118 -118 118 -32
rect 2250 1796 2486 1882
rect 2250 1732 2336 1796
rect 2400 1732 2486 1796
rect 2250 -118 2486 1732
use INV_38424460_PG0_0_0_1679678943  INV_38424460_PG0_0_0_1679678943_0
timestamp 1679679491
transform -1 0 516 0 1 0
box 0 30 516 3024
use STAGE2_INV_89403287_PG0_0_0_1679678944  STAGE2_INV_89403287_PG0_0_0_1679678944_0
timestamp 1679679491
transform -1 0 1548 0 1 0
box 0 30 1032 3024
<< labels >>
flabel metal1 s 860 588 860 588 0 FreeSerif 0 0 0 0 FOUT
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal1 s 645 1260 645 1260 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VSS
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal1 s 645 1848 645 1848 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
<< end >>
