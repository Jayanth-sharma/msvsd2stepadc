MACRO COMPARATOR
  ORIGIN 0 0 ;
  FOREIGN COMPARATOR 0 0 ;
  SIZE 19.51 BY 15.71 ;
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.6 7 17.8 7.28 ;
      LAYER M2 ;
        RECT 16.6 7.84 17.8 8.12 ;
      LAYER M2 ;
        RECT 17.04 7 17.36 7.28 ;
      LAYER M3 ;
        RECT 17.06 7.14 17.34 7.98 ;
      LAYER M2 ;
        RECT 17.04 7.84 17.36 8.12 ;
    END
  END OUT
  PIN VBIAS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
    END
  END VBIAS
  OBS 
  LAYER M2 ;
        RECT 5.42 6.58 6.62 6.86 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M2 ;
        RECT 9.72 12.04 10.92 12.32 ;
  LAYER M2 ;
        RECT 10.16 2.8 10.48 3.08 ;
  LAYER M3 ;
        RECT 10.18 2.94 10.46 12.18 ;
  LAYER M2 ;
        RECT 10.16 12.04 10.48 12.32 ;
  LAYER M2 ;
        RECT 5.86 6.58 6.18 6.86 ;
  LAYER M3 ;
        RECT 5.88 6.72 6.16 7.98 ;
  LAYER M2 ;
        RECT 5.86 7.84 6.18 8.12 ;
  LAYER M3 ;
        RECT 5.88 7.375 6.16 7.745 ;
  LAYER M2 ;
        RECT 6.02 7.42 10.32 7.7 ;
  LAYER M3 ;
        RECT 10.18 7.375 10.46 7.745 ;
  LAYER M2 ;
        RECT 5.86 6.58 6.18 6.86 ;
  LAYER M3 ;
        RECT 5.88 6.56 6.16 6.88 ;
  LAYER M2 ;
        RECT 5.86 7.84 6.18 8.12 ;
  LAYER M3 ;
        RECT 5.88 7.82 6.16 8.14 ;
  LAYER M2 ;
        RECT 5.86 6.58 6.18 6.86 ;
  LAYER M3 ;
        RECT 5.88 6.56 6.16 6.88 ;
  LAYER M2 ;
        RECT 5.86 7.84 6.18 8.12 ;
  LAYER M3 ;
        RECT 5.88 7.82 6.16 8.14 ;
  LAYER M2 ;
        RECT 5.86 6.58 6.18 6.86 ;
  LAYER M3 ;
        RECT 5.88 6.56 6.16 6.88 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 7.84 6.18 8.12 ;
  LAYER M3 ;
        RECT 5.88 7.82 6.16 8.14 ;
  LAYER M2 ;
        RECT 10.16 7.42 10.48 7.7 ;
  LAYER M3 ;
        RECT 10.18 7.4 10.46 7.72 ;
  LAYER M2 ;
        RECT 5.86 6.58 6.18 6.86 ;
  LAYER M3 ;
        RECT 5.88 6.56 6.16 6.88 ;
  LAYER M2 ;
        RECT 5.86 7.42 6.18 7.7 ;
  LAYER M3 ;
        RECT 5.88 7.4 6.16 7.72 ;
  LAYER M2 ;
        RECT 5.86 7.84 6.18 8.12 ;
  LAYER M3 ;
        RECT 5.88 7.82 6.16 8.14 ;
  LAYER M2 ;
        RECT 10.16 7.42 10.48 7.7 ;
  LAYER M3 ;
        RECT 10.18 7.4 10.46 7.72 ;
  LAYER M2 ;
        RECT 16.6 2.8 17.8 3.08 ;
  LAYER M2 ;
        RECT 16.6 12.04 17.8 12.32 ;
  LAYER M2 ;
        RECT 16.61 2.8 16.93 3.08 ;
  LAYER M3 ;
        RECT 16.63 2.94 16.91 12.18 ;
  LAYER M2 ;
        RECT 16.61 12.04 16.93 12.32 ;
  LAYER M2 ;
        RECT 13.16 7 14.36 7.28 ;
  LAYER M2 ;
        RECT 13.16 7.84 14.36 8.12 ;
  LAYER M2 ;
        RECT 13.6 7 13.92 7.28 ;
  LAYER M3 ;
        RECT 13.62 7.14 13.9 7.98 ;
  LAYER M2 ;
        RECT 13.6 7.84 13.92 8.12 ;
  LAYER M3 ;
        RECT 16.63 7.375 16.91 7.745 ;
  LAYER M2 ;
        RECT 13.76 7.42 16.77 7.7 ;
  LAYER M3 ;
        RECT 13.62 7.375 13.9 7.745 ;
  LAYER M2 ;
        RECT 13.6 7.42 13.92 7.7 ;
  LAYER M3 ;
        RECT 13.62 7.4 13.9 7.72 ;
  LAYER M2 ;
        RECT 16.61 7.42 16.93 7.7 ;
  LAYER M3 ;
        RECT 16.63 7.4 16.91 7.72 ;
  LAYER M2 ;
        RECT 13.6 7.42 13.92 7.7 ;
  LAYER M3 ;
        RECT 13.62 7.4 13.9 7.72 ;
  LAYER M2 ;
        RECT 16.61 7.42 16.93 7.7 ;
  LAYER M3 ;
        RECT 16.63 7.4 16.91 7.72 ;
  LAYER M2 ;
        RECT 1.98 7.84 3.18 8.12 ;
  LAYER M3 ;
        RECT 5.45 2.78 5.73 7.3 ;
  LAYER M2 ;
        RECT 3.01 7.84 4.73 8.12 ;
  LAYER M3 ;
        RECT 4.59 7.56 4.87 7.98 ;
  LAYER M4 ;
        RECT 4.73 7.16 5.59 7.96 ;
  LAYER M3 ;
        RECT 5.45 7.14 5.73 7.56 ;
  LAYER M2 ;
        RECT 4.57 7.84 4.89 8.12 ;
  LAYER M3 ;
        RECT 4.59 7.82 4.87 8.14 ;
  LAYER M3 ;
        RECT 4.59 7.375 4.87 7.745 ;
  LAYER M4 ;
        RECT 4.565 7.16 4.895 7.96 ;
  LAYER M3 ;
        RECT 5.45 7.375 5.73 7.745 ;
  LAYER M4 ;
        RECT 5.425 7.16 5.755 7.96 ;
  LAYER M2 ;
        RECT 4.57 7.84 4.89 8.12 ;
  LAYER M3 ;
        RECT 4.59 7.82 4.87 8.14 ;
  LAYER M3 ;
        RECT 4.59 7.375 4.87 7.745 ;
  LAYER M4 ;
        RECT 4.565 7.16 4.895 7.96 ;
  LAYER M3 ;
        RECT 5.45 7.375 5.73 7.745 ;
  LAYER M4 ;
        RECT 5.425 7.16 5.755 7.96 ;
  LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
  LAYER M2 ;
        RECT 1.55 8.26 3.61 8.54 ;
  LAYER M2 ;
        RECT 4.99 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 1.56 7 1.88 7.28 ;
  LAYER M3 ;
        RECT 1.58 7.14 1.86 8.4 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M2 ;
        RECT 3.44 8.26 5.16 8.54 ;
  LAYER M2 ;
        RECT 1.56 7 1.88 7.28 ;
  LAYER M3 ;
        RECT 1.58 6.98 1.86 7.3 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 7 1.88 7.28 ;
  LAYER M3 ;
        RECT 1.58 6.98 1.86 7.3 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 7 1.88 7.28 ;
  LAYER M3 ;
        RECT 1.58 6.98 1.86 7.3 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.56 7 1.88 7.28 ;
  LAYER M3 ;
        RECT 1.58 6.98 1.86 7.3 ;
  LAYER M2 ;
        RECT 1.56 8.26 1.88 8.54 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 8.56 ;
  LAYER M2 ;
        RECT 1.98 12.04 3.18 12.32 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M2 ;
        RECT 13.16 2.8 14.36 3.08 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 9.72 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 13.16 12.04 14.36 12.32 ;
  LAYER M2 ;
        RECT 12.04 2.8 13.33 3.08 ;
  LAYER M1 ;
        RECT 11.915 2.94 12.165 7.14 ;
  LAYER M2 ;
        RECT 10.75 7 12.04 7.28 ;
  LAYER M2 ;
        RECT 10.59 7 10.91 7.28 ;
  LAYER M3 ;
        RECT 10.61 7.14 10.89 7.98 ;
  LAYER M2 ;
        RECT 10.59 7.84 10.91 8.12 ;
  LAYER M1 ;
        RECT 11.915 7.14 12.165 12.18 ;
  LAYER M2 ;
        RECT 12.04 12.04 13.33 12.32 ;
  LAYER M1 ;
        RECT 11.915 2.855 12.165 3.025 ;
  LAYER M2 ;
        RECT 11.87 2.8 12.21 3.08 ;
  LAYER M1 ;
        RECT 11.915 7.055 12.165 7.225 ;
  LAYER M2 ;
        RECT 11.87 7 12.21 7.28 ;
  LAYER M1 ;
        RECT 11.915 2.855 12.165 3.025 ;
  LAYER M2 ;
        RECT 11.87 2.8 12.21 3.08 ;
  LAYER M1 ;
        RECT 11.915 7.055 12.165 7.225 ;
  LAYER M2 ;
        RECT 11.87 7 12.21 7.28 ;
  LAYER M1 ;
        RECT 11.915 2.855 12.165 3.025 ;
  LAYER M2 ;
        RECT 11.87 2.8 12.21 3.08 ;
  LAYER M1 ;
        RECT 11.915 7.055 12.165 7.225 ;
  LAYER M2 ;
        RECT 11.87 7 12.21 7.28 ;
  LAYER M2 ;
        RECT 10.59 7 10.91 7.28 ;
  LAYER M3 ;
        RECT 10.61 6.98 10.89 7.3 ;
  LAYER M2 ;
        RECT 10.59 7.84 10.91 8.12 ;
  LAYER M3 ;
        RECT 10.61 7.82 10.89 8.14 ;
  LAYER M1 ;
        RECT 11.915 2.855 12.165 3.025 ;
  LAYER M2 ;
        RECT 11.87 2.8 12.21 3.08 ;
  LAYER M1 ;
        RECT 11.915 7.055 12.165 7.225 ;
  LAYER M2 ;
        RECT 11.87 7 12.21 7.28 ;
  LAYER M2 ;
        RECT 10.59 7 10.91 7.28 ;
  LAYER M3 ;
        RECT 10.61 6.98 10.89 7.3 ;
  LAYER M2 ;
        RECT 10.59 7.84 10.91 8.12 ;
  LAYER M3 ;
        RECT 10.61 7.82 10.89 8.14 ;
  LAYER M1 ;
        RECT 11.915 2.855 12.165 3.025 ;
  LAYER M2 ;
        RECT 11.87 2.8 12.21 3.08 ;
  LAYER M1 ;
        RECT 11.915 7.055 12.165 7.225 ;
  LAYER M2 ;
        RECT 11.87 7 12.21 7.28 ;
  LAYER M1 ;
        RECT 11.915 12.095 12.165 12.265 ;
  LAYER M2 ;
        RECT 11.87 12.04 12.21 12.32 ;
  LAYER M2 ;
        RECT 10.59 7 10.91 7.28 ;
  LAYER M3 ;
        RECT 10.61 6.98 10.89 7.3 ;
  LAYER M2 ;
        RECT 10.59 7.84 10.91 8.12 ;
  LAYER M3 ;
        RECT 10.61 7.82 10.89 8.14 ;
  LAYER M1 ;
        RECT 11.915 2.855 12.165 3.025 ;
  LAYER M2 ;
        RECT 11.87 2.8 12.21 3.08 ;
  LAYER M1 ;
        RECT 11.915 7.055 12.165 7.225 ;
  LAYER M2 ;
        RECT 11.87 7 12.21 7.28 ;
  LAYER M1 ;
        RECT 11.915 12.095 12.165 12.265 ;
  LAYER M2 ;
        RECT 11.87 12.04 12.21 12.32 ;
  LAYER M2 ;
        RECT 10.59 7 10.91 7.28 ;
  LAYER M3 ;
        RECT 10.61 6.98 10.89 7.3 ;
  LAYER M2 ;
        RECT 10.59 7.84 10.91 8.12 ;
  LAYER M3 ;
        RECT 10.61 7.82 10.89 8.14 ;
  LAYER M1 ;
        RECT 10.625 3.695 10.875 7.225 ;
  LAYER M1 ;
        RECT 10.625 2.435 10.875 3.445 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 10.195 3.695 10.445 7.225 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.765 2.435 10.015 3.445 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 9.29 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 9.72 0.7 10.92 0.98 ;
  LAYER M2 ;
        RECT 9.72 7 10.92 7.28 ;
  LAYER M2 ;
        RECT 9.72 2.8 10.92 3.08 ;
  LAYER M3 ;
        RECT 9.75 0.68 10.03 6.88 ;
  LAYER M1 ;
        RECT 14.065 3.695 14.315 7.225 ;
  LAYER M1 ;
        RECT 14.065 2.435 14.315 3.445 ;
  LAYER M1 ;
        RECT 14.065 0.335 14.315 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M2 ;
        RECT 12.73 6.58 14.79 6.86 ;
  LAYER M2 ;
        RECT 13.16 0.7 14.36 0.98 ;
  LAYER M2 ;
        RECT 13.16 7 14.36 7.28 ;
  LAYER M2 ;
        RECT 13.16 2.8 14.36 3.08 ;
  LAYER M3 ;
        RECT 13.19 0.68 13.47 6.88 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 9.765 7.895 10.015 11.425 ;
  LAYER M1 ;
        RECT 9.765 11.675 10.015 12.685 ;
  LAYER M1 ;
        RECT 9.765 13.775 10.015 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M2 ;
        RECT 9.29 8.26 11.35 8.54 ;
  LAYER M2 ;
        RECT 9.72 14.14 10.92 14.42 ;
  LAYER M2 ;
        RECT 9.72 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 9.72 12.04 10.92 12.32 ;
  LAYER M3 ;
        RECT 9.75 8.24 10.03 14.44 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 11.425 ;
  LAYER M1 ;
        RECT 14.065 11.675 14.315 12.685 ;
  LAYER M1 ;
        RECT 14.065 13.775 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.495 7.895 14.745 11.425 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 11.425 ;
  LAYER M1 ;
        RECT 13.205 11.675 13.455 12.685 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 14.785 ;
  LAYER M1 ;
        RECT 12.775 7.895 13.025 11.425 ;
  LAYER M2 ;
        RECT 12.73 8.26 14.79 8.54 ;
  LAYER M2 ;
        RECT 13.16 14.14 14.36 14.42 ;
  LAYER M2 ;
        RECT 13.16 7.84 14.36 8.12 ;
  LAYER M2 ;
        RECT 13.16 12.04 14.36 12.32 ;
  LAYER M3 ;
        RECT 13.19 8.24 13.47 14.44 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 5.465 3.695 5.715 7.225 ;
  LAYER M1 ;
        RECT 5.465 2.435 5.715 3.445 ;
  LAYER M1 ;
        RECT 5.465 0.335 5.715 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 4.56 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 4.13 6.16 7.91 6.44 ;
  LAYER M2 ;
        RECT 4.56 0.7 7.48 0.98 ;
  LAYER M3 ;
        RECT 5.45 2.78 5.73 7.3 ;
  LAYER M2 ;
        RECT 5.42 6.58 6.62 6.86 ;
  LAYER M3 ;
        RECT 6.31 0.68 6.59 6.46 ;
  LAYER M1 ;
        RECT 16.645 3.695 16.895 7.225 ;
  LAYER M1 ;
        RECT 16.645 2.435 16.895 3.445 ;
  LAYER M1 ;
        RECT 16.645 0.335 16.895 1.345 ;
  LAYER M1 ;
        RECT 16.215 3.695 16.465 7.225 ;
  LAYER M1 ;
        RECT 17.075 3.695 17.325 7.225 ;
  LAYER M1 ;
        RECT 17.505 3.695 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.505 2.435 17.755 3.445 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 1.345 ;
  LAYER M1 ;
        RECT 17.935 3.695 18.185 7.225 ;
  LAYER M2 ;
        RECT 16.17 6.58 18.23 6.86 ;
  LAYER M2 ;
        RECT 16.6 0.7 17.8 0.98 ;
  LAYER M2 ;
        RECT 16.6 7 17.8 7.28 ;
  LAYER M2 ;
        RECT 16.6 2.8 17.8 3.08 ;
  LAYER M3 ;
        RECT 17.49 0.68 17.77 6.88 ;
  LAYER M1 ;
        RECT 16.645 7.895 16.895 11.425 ;
  LAYER M1 ;
        RECT 16.645 11.675 16.895 12.685 ;
  LAYER M1 ;
        RECT 16.645 13.775 16.895 14.785 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M1 ;
        RECT 17.075 7.895 17.325 11.425 ;
  LAYER M1 ;
        RECT 17.505 7.895 17.755 11.425 ;
  LAYER M1 ;
        RECT 17.505 11.675 17.755 12.685 ;
  LAYER M1 ;
        RECT 17.505 13.775 17.755 14.785 ;
  LAYER M1 ;
        RECT 17.935 7.895 18.185 11.425 ;
  LAYER M2 ;
        RECT 16.17 8.26 18.23 8.54 ;
  LAYER M2 ;
        RECT 16.6 14.14 17.8 14.42 ;
  LAYER M2 ;
        RECT 16.6 7.84 17.8 8.12 ;
  LAYER M2 ;
        RECT 16.6 12.04 17.8 12.32 ;
  LAYER M3 ;
        RECT 17.49 8.24 17.77 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 2.75 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.7 2.32 0.98 ;
  LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M3 ;
        RECT 2.01 0.68 2.29 6.88 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M2 ;
        RECT 1.98 14.14 3.18 14.42 ;
  LAYER M2 ;
        RECT 1.98 7.84 3.18 8.12 ;
  LAYER M2 ;
        RECT 1.98 12.04 3.18 12.32 ;
  LAYER M2 ;
        RECT 1.55 8.26 3.61 8.54 ;
  LAYER M1 ;
        RECT 5.465 7.895 5.715 11.425 ;
  LAYER M1 ;
        RECT 5.465 11.675 5.715 12.685 ;
  LAYER M1 ;
        RECT 5.465 13.775 5.715 14.785 ;
  LAYER M1 ;
        RECT 5.035 7.895 5.285 11.425 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M2 ;
        RECT 5.42 14.14 6.62 14.42 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M2 ;
        RECT 4.99 8.26 7.05 8.54 ;
  END 
END COMPARATOR
