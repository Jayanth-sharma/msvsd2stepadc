magic
tech sky130A
magscale 1 2
timestamp 1678040207
<< pwell >>
rect 478 436 532 444
rect 478 356 540 436
<< locali >>
rect 474 448 1536 458
rect 474 434 1468 448
rect 474 370 484 434
rect 536 388 1468 434
rect 536 370 1536 388
rect 474 360 1536 370
<< viali >>
rect 484 370 536 434
rect 1468 388 1536 448
<< metal1 >>
rect 310 1136 1568 1206
rect 354 1048 1568 1136
rect 354 902 406 1048
rect 496 1000 554 1002
rect 496 948 556 1000
rect 498 946 556 948
rect 354 836 502 902
rect 762 898 796 1048
rect 900 950 964 1004
rect 1170 912 1210 1048
rect 1318 952 1382 1006
rect 762 810 910 898
rect 1170 816 1336 912
rect 1462 800 1522 804
rect 556 722 700 794
rect 958 788 1102 794
rect 958 722 1108 788
rect 1380 728 1528 800
rect 464 626 558 680
rect 464 434 546 626
rect 464 370 484 434
rect 536 370 546 434
rect 464 162 546 370
rect 638 448 698 722
rect 898 670 962 676
rect 884 622 962 670
rect 884 448 958 622
rect 638 366 958 448
rect 638 122 698 366
rect 884 166 958 366
rect 1048 458 1108 722
rect 1314 676 1388 678
rect 1314 622 1392 676
rect 1314 458 1388 622
rect 1048 376 1388 458
rect 526 50 698 122
rect 1048 116 1108 376
rect 1314 174 1388 376
rect 1462 464 1522 728
rect 1462 448 1600 464
rect 1462 388 1468 448
rect 1536 388 1600 448
rect 1462 376 1600 388
rect 1314 170 1378 174
rect 1462 132 1522 376
rect 950 44 1108 116
rect 1368 60 1522 132
rect 318 34 468 38
rect 314 -50 468 34
rect 748 -24 898 34
rect 314 -194 354 -50
rect 744 -54 898 -24
rect 1170 -54 1320 34
rect 468 -150 532 -96
rect 744 -194 784 -54
rect 888 -146 952 -92
rect 1170 -194 1210 -54
rect 1314 -142 1378 -88
rect 278 -360 1564 -194
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1678040207
transform 1 0 921 0 1 36
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1678040207
transform 1 0 527 0 1 813
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM3
timestamp 1678040207
transform 1 0 1345 0 1 40
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM4
timestamp 1678040207
transform 1 0 933 0 1 815
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 1678040207
transform 1 0 497 0 1 32
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM6
timestamp 1678040207
transform 1 0 1353 0 1 815
box -211 -319 211 319
<< labels >>
rlabel space 1530 1072 1570 1202 3 vdd
port 1 e
rlabel space 1560 370 1598 468 3 out
port 2 e
rlabel space 1520 -368 1564 -188 3 vss
port 3 e
<< end >>
