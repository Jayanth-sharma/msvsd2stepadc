* SPICE3 file created from TWOBIT_DAC_0.ext - technology: sky130A
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.subckt Twobit_DAC OUT VDD GND X1_INP1 X1_INP2 X2_INP1 X2_INP2 D0 D1
X0 SWITCH_PG0_0_0_1680779960_0/m1_226_2912# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# m1_2322_1568# VDD sky130_fd_pr__pfet_01v8 ad=6.678e+11p pd=6.1e+06u as=1.3734e+12p ps=1.226e+07u w=1.26e+06u l=150000u
X1 m1_2322_1568# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_226_2912# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X2 m1_2322_1568# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_656_2912# GND sky130_fd_pr__nfet_01v8 ad=8.442e+11p pd=8.98e+06u as=3.339e+11p ps=3.58e+06u w=630000u l=150000u
X3 SWITCH_PG0_0_0_1680779960_0/m1_656_2912# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# m1_2322_1568# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X4 SWITCH_PG0_0_0_1680779960_0/m1_226_2912# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# m1_2322_1568# GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=0p ps=0u w=630000u l=150000u
X5 m1_2322_1568# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# SWITCH_PG0_0_0_1680779960_0/m1_226_2912# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X6 SWITCH_PG0_0_0_1680779960_0/m1_774_2072# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# GND GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=2.0034e+12p ps=2.148e+07u w=630000u l=150000u
X7 GND SWITCH_PG0_0_0_1680779960_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X8 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# D0 GND GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=0p ps=0u w=630000u l=150000u
X9 GND D0 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X10 VDD D0 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# VDD sky130_fd_pr__pfet_01v8 ad=4.0068e+12p pd=3.66e+07u as=3.528e+11p ps=3.08e+06u w=1.26e+06u l=150000u
X11 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# D0 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X12 VDD SWITCH_PG0_0_0_1680779960_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.528e+11p ps=3.08e+06u w=1.26e+06u l=150000u
X13 SWITCH_PG0_0_0_1680779960_0/m1_774_2072# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X14 m1_2322_1568# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# SWITCH_PG0_0_0_1680779960_0/m1_656_2912# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.528e+11p ps=3.08e+06u w=1.26e+06u l=150000u
X15 SWITCH_PG0_0_0_1680779960_0/m1_656_2912# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# m1_2322_1568# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X16 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# GND GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=0p ps=0u w=630000u l=150000u
X17 GND SWITCH_PG0_1_0_1680779961_0/m1_430_3920# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X18 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# D0 GND GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=0p ps=0u w=630000u l=150000u
X19 GND D0 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X20 VDD SWITCH_PG0_1_0_1680779961_0/m1_430_3920# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.528e+11p ps=3.08e+06u w=1.26e+06u l=150000u
X21 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X22 VDD D0 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.528e+11p ps=3.08e+06u w=1.26e+06u l=150000u
X23 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# D0 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X24 m1_1376_1652# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# SWITCH_PG0_1_0_1680779961_0/li_577_2923# VDD sky130_fd_pr__pfet_01v8 ad=1.6884e+12p pd=1.528e+07u as=3.528e+11p ps=3.08e+06u w=1.26e+06u l=150000u
X25 SWITCH_PG0_1_0_1680779961_0/li_577_2923# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# m1_1376_1652# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X26 SWITCH_PG0_1_0_1680779961_0/m1_312_2912# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# m1_1376_1652# VDD sky130_fd_pr__pfet_01v8 ad=6.678e+11p pd=6.1e+06u as=0p ps=0u w=1.26e+06u l=150000u
X27 m1_1376_1652# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# SWITCH_PG0_1_0_1680779961_0/m1_312_2912# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X28 m1_1376_1652# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# SWITCH_PG0_1_0_1680779961_0/li_577_2923# GND sky130_fd_pr__nfet_01v8 ad=6.867e+11p pd=7.22e+06u as=3.339e+11p ps=3.58e+06u w=630000u l=150000u
X29 SWITCH_PG0_1_0_1680779961_0/li_577_2923# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# m1_1376_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X30 SWITCH_PG0_1_0_1680779961_0/m1_312_2912# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# m1_1376_1652# GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=0p ps=0u w=630000u l=150000u
X31 m1_1376_1652# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# SWITCH_PG0_1_0_1680779961_0/m1_312_2912# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X32 OUT SWITCH_PG0_2_0_1680779962_0/m1_430_3920# m1_2322_1568# GND sky130_fd_pr__nfet_01v8 ad=5.103e+11p pd=5.4e+06u as=0p ps=0u w=630000u l=150000u
X33 m1_2322_1568# SWITCH_PG0_2_0_1680779962_0/m1_430_3920# OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X34 m1_1376_1652# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X35 OUT SWITCH_PG0_2_0_1680779962_0/m1_774_2072# m1_1376_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X36 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# SWITCH_PG0_2_0_1680779962_0/m1_430_3920# GND GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=0p ps=0u w=630000u l=150000u
X37 GND SWITCH_PG0_2_0_1680779962_0/m1_430_3920# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X38 m1_1376_1652# SWITCH_PG0_2_0_1680779962_0/m1_430_3920# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.0206e+12p ps=9.18e+06u w=1.26e+06u l=150000u
X39 OUT SWITCH_PG0_2_0_1680779962_0/m1_430_3920# m1_1376_1652# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X40 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# D1 GND GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=0p ps=0u w=630000u l=150000u
X41 GND D1 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X42 VDD SWITCH_PG0_2_0_1680779962_0/m1_430_3920# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.528e+11p ps=3.08e+06u w=1.26e+06u l=150000u
X43 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# SWITCH_PG0_2_0_1680779962_0/m1_430_3920# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X44 VDD D1 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.528e+11p ps=3.08e+06u w=1.26e+06u l=150000u
X45 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# D1 VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X46 OUT SWITCH_PG0_2_0_1680779962_0/m1_774_2072# m1_2322_1568# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X47 m1_2322_1568# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# OUT VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
C0 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# VDD 4.31fF
C1 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# 0.00fF
C2 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# D1 0.00fF
C3 VDD OUT 0.74fF
C4 VDD SWITCH_PG0_0_0_1680779960_0/m1_226_2912# 0.25fF
C5 m1_2322_1568# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 0.29fF
C6 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# OUT 0.00fF
C7 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# VDD 1.93fF
C8 m1_1376_1652# X2_INP1 0.00fF
C9 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 0.01fF
C10 X2_INP1 m1_2322_1568# 0.04fF
C11 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# 0.03fF
C12 X2_INP1 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.00fF
C13 SWITCH_PG0_1_0_1680779961_0/m1_312_2912# VDD 0.27fF
C14 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# OUT 0.00fF
C15 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_226_2912# 0.11fF
C16 SWITCH_PG0_1_0_1680779961_0/m1_312_2912# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# 0.11fF
C17 VDD SWITCH_PG0_0_0_1680779960_0/m1_430_3920# 4.07fF
C18 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# D0 0.08fF
C19 VDD D0 3.87fF
C20 X2_INP2 SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 0.00fF
C21 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# D0 0.00fF
C22 SWITCH_PG0_0_0_1680779960_0/m1_656_2912# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 0.11fF
C23 SWITCH_PG0_1_0_1680779961_0/li_577_2923# VDD 0.30fF
C24 m1_1376_1652# SWITCH_PG0_2_0_1680779962_0/m1_430_3920# 0.10fF
C25 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# SWITCH_PG0_1_0_1680779961_0/li_577_2923# 0.10fF
C26 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# X1_INP1 0.00fF
C27 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# m1_2322_1568# 0.56fF
C28 D0 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# 0.25fF
C29 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.40fF
C30 m1_1376_1652# OUT 1.80fF
C31 X1_INP1 OUT 0.00fF
C32 m1_2322_1568# OUT 1.55fF
C33 SWITCH_PG0_1_0_1680779961_0/m1_312_2912# SWITCH_PG0_1_0_1680779961_0/li_577_2923# 0.09fF
C34 m1_2322_1568# SWITCH_PG0_0_0_1680779960_0/m1_226_2912# 1.72fF
C35 m1_1376_1652# VDD 1.17fF
C36 VDD X1_INP1 0.06fF
C37 m1_2322_1568# VDD 2.34fF
C38 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# OUT 0.29fF
C39 m1_1376_1652# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# 0.23fF
C40 VDD SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 1.96fF
C41 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# m1_2322_1568# 0.00fF
C42 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# X1_INP2 0.00fF
C43 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.04fF
C44 m1_1376_1652# SWITCH_PG0_1_0_1680779961_0/m1_312_2912# 1.61fF
C45 X1_INP2 OUT 0.00fF
C46 m1_1376_1652# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# 0.00fF
C47 VDD X1_INP2 0.01fF
C48 m1_2322_1568# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# 0.36fF
C49 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# D1 0.20fF
C50 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# 0.04fF
C51 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# SWITCH_PG0_0_0_1680779960_0/m1_430_3920# 0.00fF
C52 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# X2_INP2 0.00fF
C53 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# OUT 0.00fF
C54 D1 VDD 0.82fF
C55 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# VDD 3.84fF
C56 X2_INP2 OUT 0.00fF
C57 VDD X2_INP2 0.04fF
C58 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# SWITCH_PG0_1_0_1680779961_0/m1_774_2072# 0.49fF
C59 SWITCH_PG0_0_0_1680779960_0/m1_656_2912# SWITCH_PG0_0_0_1680779960_0/m1_226_2912# 0.08fF
C60 D0 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.00fF
C61 VDD SWITCH_PG0_0_0_1680779960_0/m1_656_2912# 0.30fF
C62 m1_1376_1652# SWITCH_PG0_1_0_1680779961_0/li_577_2923# 1.67fF
C63 SWITCH_PG0_1_0_1680779961_0/m1_312_2912# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# 0.11fF
C64 D1 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# 0.00fF
C65 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 0.01fF
C66 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# X2_INP2 0.01fF
C67 m1_1376_1652# X1_INP1 0.06fF
C68 m1_1376_1652# m1_2322_1568# 0.07fF
C69 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_656_2912# 0.35fF
C70 m1_2322_1568# X1_INP1 0.00fF
C71 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# X2_INP1 0.02fF
C72 SWITCH_PG0_0_0_1680779960_0/m1_774_2072# OUT 0.00fF
C73 SWITCH_PG0_0_0_1680779960_0/m1_226_2912# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 0.11fF
C74 m1_1376_1652# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.11fF
C75 D1 D0 0.78fF
C76 X1_INP1 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.00fF
C77 m1_2322_1568# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.18fF
C78 VDD SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 1.92fF
C79 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# D0 0.23fF
C80 X2_INP1 OUT 0.00fF
C81 X2_INP1 VDD 0.21fF
C82 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# SWITCH_PG0_1_0_1680779961_0/li_577_2923# 0.36fF
C83 m1_2322_1568# X1_INP2 0.00fF
C84 X1_INP2 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.00fF
C85 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 0.40fF
C86 m1_1376_1652# SWITCH_PG0_1_0_1680779961_0/m1_430_3920# 0.36fF
C87 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# m1_2322_1568# 0.00fF
C88 D1 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.00fF
C89 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# SWITCH_PG0_2_0_1680779962_0/m1_774_2072# 0.00fF
C90 m1_2322_1568# SWITCH_PG0_0_0_1680779960_0/m1_656_2912# 1.62fF
C91 D0 SWITCH_PG0_0_0_1680779960_0/m1_774_2072# 0.00fF
C92 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# X2_INP2 0.00fF
C93 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# OUT 0.36fF
C94 X1_INP2 GND 0.24fF
C95 X1_INP1 GND 0.17fF
C96 X2_INP2 GND 0.34fF
C97 X2_INP1 GND 0.14fF
C98 SWITCH_PG0_2_0_1680779962_0/m1_774_2072# GND 1.37fF
C99 OUT GND 0.11fF
C100 D1 GND 0.71fF
C101 VDD GND 41.82fF
C102 SWITCH_PG0_2_0_1680779962_0/m1_430_3920# GND 1.76fF
C103 SWITCH_PG0_1_0_1680779961_0/m1_774_2072# GND 1.26fF
C104 SWITCH_PG0_1_0_1680779961_0/m1_312_2912# GND 0.08fF
C105 SWITCH_PG0_1_0_1680779961_0/li_577_2923# GND 0.05fF
C106 SWITCH_PG0_1_0_1680779961_0/m1_430_3920# GND 1.97fF
C107 SWITCH_PG0_0_0_1680779960_0/m1_774_2072# GND 1.52fF
C108 SWITCH_PG0_0_0_1680779960_0/m1_656_2912# GND 0.02fF
C109 SWITCH_PG0_0_0_1680779960_0/m1_430_3920# GND 1.83fF
C110 SWITCH_PG0_0_0_1680779960_0/m1_226_2912# GND 0.10fF
.ends  Twobit_DAC

x1 OUT VDD GND X1_INP1 X1_INP2 X2_INP1 X2_INP2 D0 D1 Twobit_DAC 
V1 X2_INP2 GND 0.1
V2 X1_INP1 GND 2.47
V3 X1_INP2 GND 1.57
V4 X2_INP1 GND 0.75
V5 D0 GND pulse(0 1.8 0n 1p 1p 5u 10u)
V6 VDD GND 3.3
V7 D1 GND pulse(0 1.8 0n 1p 1p 10u 20u)

.tran 1n 20u
.control
run
plot v(D0) v(D1) v(OUT)
.endc

