MACRO TWO_BIT_RES_DAC
  ORIGIN 0 0 ;
  FOREIGN TWO_BIT_RES_DAC 0 0 ;
  SIZE 19.51 BY 45.95 ;
  PIN D0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 27.16 2.32 27.44 ;
      LAYER M2 ;
        RECT 2.84 27.16 4.04 27.44 ;
      LAYER M2 ;
        RECT 2.15 27.16 3.01 27.44 ;
      LAYER M2 ;
        RECT 1.12 42.28 2.32 42.56 ;
      LAYER M2 ;
        RECT 2.84 42.28 4.04 42.56 ;
      LAYER M2 ;
        RECT 2.15 42.28 3.01 42.56 ;
      LAYER M2 ;
        RECT 2.42 27.16 2.74 27.44 ;
      LAYER M3 ;
        RECT 2.44 27.3 2.72 42.42 ;
      LAYER M2 ;
        RECT 2.42 42.28 2.74 42.56 ;
    END
  END D0
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
      LAYER M2 ;
        RECT 2.84 2.8 4.04 3.08 ;
      LAYER M2 ;
        RECT 2.15 2.8 3.01 3.08 ;
    END
  END D1
  PIN OUT_V
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
      LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
      LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
      LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
      LAYER M2 ;
        RECT 8.44 7 8.76 7.28 ;
      LAYER M3 ;
        RECT 8.46 7.14 8.74 7.98 ;
      LAYER M2 ;
        RECT 8.44 7.84 8.76 8.12 ;
      LAYER M3 ;
        RECT 4.16 8.635 4.44 9.005 ;
      LAYER M2 ;
        RECT 4.3 8.68 6.02 8.96 ;
      LAYER M3 ;
        RECT 5.88 8.635 6.16 9.005 ;
      LAYER M2 ;
        RECT 6.02 8.68 8.17 8.96 ;
      LAYER M3 ;
        RECT 8.03 7.98 8.31 8.82 ;
      LAYER M2 ;
        RECT 8.01 7.84 8.33 8.12 ;
    END
  END OUT_V
  OBS 
  LAYER M3 ;
        RECT 4.16 38.48 4.44 44.68 ;
  LAYER M3 ;
        RECT 5.88 38.48 6.16 44.68 ;
  LAYER M3 ;
        RECT 4.16 41.395 4.44 41.765 ;
  LAYER M2 ;
        RECT 4.3 41.44 6.02 41.72 ;
  LAYER M3 ;
        RECT 5.88 41.395 6.16 41.765 ;
  LAYER M4 ;
        RECT 10.585 43.7 18.225 44.5 ;
  LAYER M3 ;
        RECT 5.88 43.915 6.16 44.285 ;
  LAYER M4 ;
        RECT 6.02 43.7 10.75 44.5 ;
  LAYER M3 ;
        RECT 5.88 43.915 6.16 44.285 ;
  LAYER M4 ;
        RECT 5.855 43.7 6.185 44.5 ;
  LAYER M3 ;
        RECT 5.88 43.915 6.16 44.285 ;
  LAYER M4 ;
        RECT 5.855 43.7 6.185 44.5 ;
  LAYER M2 ;
        RECT 6.28 30.52 7.48 30.8 ;
  LAYER M3 ;
        RECT 9.32 30.92 9.6 37.12 ;
  LAYER M2 ;
        RECT 7.31 30.52 9.46 30.8 ;
  LAYER M3 ;
        RECT 9.32 30.66 9.6 31.08 ;
  LAYER M4 ;
        RECT 10.585 32.36 18.225 33.16 ;
  LAYER M4 ;
        RECT 10.585 34.88 18.225 35.68 ;
  LAYER M4 ;
        RECT 14.025 32.36 14.355 33.16 ;
  LAYER M3 ;
        RECT 14.05 32.76 14.33 35.28 ;
  LAYER M4 ;
        RECT 14.025 34.88 14.355 35.68 ;
  LAYER M3 ;
        RECT 9.32 32.575 9.6 32.945 ;
  LAYER M4 ;
        RECT 9.46 32.36 10.75 33.16 ;
  LAYER M3 ;
        RECT 9.32 32.575 9.6 32.945 ;
  LAYER M4 ;
        RECT 9.295 32.36 9.625 33.16 ;
  LAYER M3 ;
        RECT 9.32 32.575 9.6 32.945 ;
  LAYER M4 ;
        RECT 9.295 32.36 9.625 33.16 ;
  LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 6.88 ;
  LAYER M3 ;
        RECT 4.16 3.595 4.44 3.965 ;
  LAYER M2 ;
        RECT 4.3 3.64 6.02 3.92 ;
  LAYER M3 ;
        RECT 5.88 3.595 6.16 3.965 ;
  LAYER M3 ;
        RECT 4.16 30.92 4.44 37.12 ;
  LAYER M3 ;
        RECT 5.88 30.92 6.16 37.12 ;
  LAYER M2 ;
        RECT 8 37.24 9.2 37.52 ;
  LAYER M2 ;
        RECT 8 38.08 9.2 38.36 ;
  LAYER M2 ;
        RECT 8.44 37.24 8.76 37.52 ;
  LAYER M3 ;
        RECT 8.46 37.38 8.74 38.22 ;
  LAYER M2 ;
        RECT 8.44 38.08 8.76 38.36 ;
  LAYER M3 ;
        RECT 4.16 36.355 4.44 36.725 ;
  LAYER M2 ;
        RECT 4.3 36.4 6.02 36.68 ;
  LAYER M3 ;
        RECT 5.88 36.355 6.16 36.725 ;
  LAYER M2 ;
        RECT 6.02 36.4 8.17 36.68 ;
  LAYER M3 ;
        RECT 8.03 36.54 8.31 37.38 ;
  LAYER M2 ;
        RECT 8.01 37.24 8.33 37.52 ;
  LAYER M3 ;
        RECT 5.88 6.72 6.16 7.56 ;
  LAYER M4 ;
        RECT 5.59 7.16 6.02 7.96 ;
  LAYER M3 ;
        RECT 5.45 7.56 5.73 30.24 ;
  LAYER M2 ;
        RECT 5.59 30.1 6.02 30.38 ;
  LAYER M3 ;
        RECT 5.88 30.24 6.16 31.08 ;
  LAYER M2 ;
        RECT 5.43 30.1 5.75 30.38 ;
  LAYER M3 ;
        RECT 5.45 30.08 5.73 30.4 ;
  LAYER M2 ;
        RECT 5.86 30.1 6.18 30.38 ;
  LAYER M3 ;
        RECT 5.88 30.08 6.16 30.4 ;
  LAYER M3 ;
        RECT 5.45 7.375 5.73 7.745 ;
  LAYER M4 ;
        RECT 5.425 7.16 5.755 7.96 ;
  LAYER M3 ;
        RECT 5.88 7.375 6.16 7.745 ;
  LAYER M4 ;
        RECT 5.855 7.16 6.185 7.96 ;
  LAYER M2 ;
        RECT 5.43 30.1 5.75 30.38 ;
  LAYER M3 ;
        RECT 5.45 30.08 5.73 30.4 ;
  LAYER M2 ;
        RECT 5.86 30.1 6.18 30.38 ;
  LAYER M3 ;
        RECT 5.88 30.08 6.16 30.4 ;
  LAYER M3 ;
        RECT 5.45 7.375 5.73 7.745 ;
  LAYER M4 ;
        RECT 5.425 7.16 5.755 7.96 ;
  LAYER M3 ;
        RECT 5.88 7.375 6.16 7.745 ;
  LAYER M4 ;
        RECT 5.855 7.16 6.185 7.96 ;
  LAYER M3 ;
        RECT 4.16 23.36 4.44 29.56 ;
  LAYER M3 ;
        RECT 5.88 23.36 6.16 29.56 ;
  LAYER M3 ;
        RECT 4.16 26.275 4.44 26.645 ;
  LAYER M2 ;
        RECT 4.3 26.32 6.02 26.6 ;
  LAYER M3 ;
        RECT 5.88 26.275 6.16 26.645 ;
  LAYER M4 ;
        RECT 10.585 23.54 18.225 24.34 ;
  LAYER M4 ;
        RECT 10.585 21.02 18.225 21.82 ;
  LAYER M3 ;
        RECT 5.88 23.755 6.16 24.125 ;
  LAYER M4 ;
        RECT 6.02 23.54 10.75 24.34 ;
  LAYER M4 ;
        RECT 10.585 23.54 10.915 24.34 ;
  LAYER M3 ;
        RECT 10.61 21.42 10.89 23.94 ;
  LAYER M4 ;
        RECT 10.585 21.02 10.915 21.82 ;
  LAYER M3 ;
        RECT 5.88 23.755 6.16 24.125 ;
  LAYER M4 ;
        RECT 5.855 23.54 6.185 24.34 ;
  LAYER M3 ;
        RECT 5.88 23.755 6.16 24.125 ;
  LAYER M4 ;
        RECT 5.855 23.54 6.185 24.34 ;
  LAYER M3 ;
        RECT 5.88 23.755 6.16 24.125 ;
  LAYER M4 ;
        RECT 5.855 23.54 6.185 24.34 ;
  LAYER M3 ;
        RECT 10.61 21.235 10.89 21.605 ;
  LAYER M4 ;
        RECT 10.585 21.02 10.915 21.82 ;
  LAYER M3 ;
        RECT 10.61 23.755 10.89 24.125 ;
  LAYER M4 ;
        RECT 10.585 23.54 10.915 24.34 ;
  LAYER M3 ;
        RECT 5.88 23.755 6.16 24.125 ;
  LAYER M4 ;
        RECT 5.855 23.54 6.185 24.34 ;
  LAYER M3 ;
        RECT 10.61 21.235 10.89 21.605 ;
  LAYER M4 ;
        RECT 10.585 21.02 10.915 21.82 ;
  LAYER M3 ;
        RECT 10.61 23.755 10.89 24.125 ;
  LAYER M4 ;
        RECT 10.585 23.54 10.915 24.34 ;
  LAYER M2 ;
        RECT 6.28 15.4 7.48 15.68 ;
  LAYER M3 ;
        RECT 9.32 15.8 9.6 22 ;
  LAYER M2 ;
        RECT 7.31 15.4 9.46 15.68 ;
  LAYER M3 ;
        RECT 9.32 15.54 9.6 15.96 ;
  LAYER M4 ;
        RECT 10.585 9.68 18.225 10.48 ;
  LAYER M4 ;
        RECT 10.585 12.2 18.225 13 ;
  LAYER M4 ;
        RECT 14.025 9.68 14.355 10.48 ;
  LAYER M3 ;
        RECT 14.05 10.08 14.33 12.6 ;
  LAYER M4 ;
        RECT 14.025 12.2 14.355 13 ;
  LAYER M2 ;
        RECT 9.46 15.4 10.75 15.68 ;
  LAYER M3 ;
        RECT 10.61 12.6 10.89 15.54 ;
  LAYER M4 ;
        RECT 10.585 12.2 10.915 13 ;
  LAYER M2 ;
        RECT 10.59 15.4 10.91 15.68 ;
  LAYER M3 ;
        RECT 10.61 15.38 10.89 15.7 ;
  LAYER M3 ;
        RECT 10.61 12.415 10.89 12.785 ;
  LAYER M4 ;
        RECT 10.585 12.2 10.915 13 ;
  LAYER M2 ;
        RECT 10.59 15.4 10.91 15.68 ;
  LAYER M3 ;
        RECT 10.61 15.38 10.89 15.7 ;
  LAYER M3 ;
        RECT 10.61 12.415 10.89 12.785 ;
  LAYER M4 ;
        RECT 10.585 12.2 10.915 13 ;
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M3 ;
        RECT 9.32 14.28 9.6 14.7 ;
  LAYER M2 ;
        RECT 7.31 14.56 9.46 14.84 ;
  LAYER M3 ;
        RECT 4.16 15.8 4.44 22 ;
  LAYER M3 ;
        RECT 5.88 15.8 6.16 22 ;
  LAYER M2 ;
        RECT 8 22.12 9.2 22.4 ;
  LAYER M2 ;
        RECT 8 22.96 9.2 23.24 ;
  LAYER M2 ;
        RECT 8.44 22.12 8.76 22.4 ;
  LAYER M3 ;
        RECT 8.46 22.26 8.74 23.1 ;
  LAYER M2 ;
        RECT 8.44 22.96 8.76 23.24 ;
  LAYER M3 ;
        RECT 4.16 21.235 4.44 21.605 ;
  LAYER M2 ;
        RECT 4.3 21.28 6.02 21.56 ;
  LAYER M3 ;
        RECT 5.88 21.235 6.16 21.605 ;
  LAYER M2 ;
        RECT 6.02 21.28 8.17 21.56 ;
  LAYER M3 ;
        RECT 8.03 21.42 8.31 22.26 ;
  LAYER M2 ;
        RECT 8.01 22.12 8.33 22.4 ;
  LAYER M2 ;
        RECT 6.29 14.56 6.61 14.84 ;
  LAYER M3 ;
        RECT 6.31 14.7 6.59 15.12 ;
  LAYER M2 ;
        RECT 6.02 14.98 6.45 15.26 ;
  LAYER M3 ;
        RECT 5.88 15.12 6.16 15.96 ;
  LAYER M2 ;
        RECT 5.86 14.98 6.18 15.26 ;
  LAYER M3 ;
        RECT 5.88 14.96 6.16 15.28 ;
  LAYER M2 ;
        RECT 6.29 14.56 6.61 14.84 ;
  LAYER M3 ;
        RECT 6.31 14.54 6.59 14.86 ;
  LAYER M2 ;
        RECT 6.29 14.98 6.61 15.26 ;
  LAYER M3 ;
        RECT 6.31 14.96 6.59 15.28 ;
  LAYER M2 ;
        RECT 5.86 14.98 6.18 15.26 ;
  LAYER M3 ;
        RECT 5.88 14.96 6.16 15.28 ;
  LAYER M2 ;
        RECT 6.29 14.56 6.61 14.84 ;
  LAYER M3 ;
        RECT 6.31 14.54 6.59 14.86 ;
  LAYER M2 ;
        RECT 6.29 14.98 6.61 15.26 ;
  LAYER M3 ;
        RECT 6.31 14.96 6.59 15.28 ;
  LAYER M4 ;
        RECT 10.585 0.86 18.225 1.66 ;
  LAYER M2 ;
        RECT 1.12 37.24 2.32 37.52 ;
  LAYER M2 ;
        RECT 6.28 38.08 7.48 38.36 ;
  LAYER M2 ;
        RECT 8 33.04 9.2 33.32 ;
  LAYER M2 ;
        RECT 8 42.28 9.2 42.56 ;
  LAYER M2 ;
        RECT 8.01 33.04 8.33 33.32 ;
  LAYER M1 ;
        RECT 8.045 33.18 8.295 42.42 ;
  LAYER M2 ;
        RECT 8.01 42.28 8.33 42.56 ;
  LAYER M2 ;
        RECT 1.99 37.24 2.31 37.52 ;
  LAYER M1 ;
        RECT 2.025 37.38 2.275 37.8 ;
  LAYER M2 ;
        RECT 2.15 37.66 6.45 37.94 ;
  LAYER M3 ;
        RECT 6.31 37.8 6.59 38.22 ;
  LAYER M2 ;
        RECT 6.29 38.08 6.61 38.36 ;
  LAYER M2 ;
        RECT 6.45 37.66 8.17 37.94 ;
  LAYER M1 ;
        RECT 8.045 37.715 8.295 37.885 ;
  LAYER M1 ;
        RECT 2.025 37.295 2.275 37.465 ;
  LAYER M2 ;
        RECT 1.98 37.24 2.32 37.52 ;
  LAYER M1 ;
        RECT 2.025 37.715 2.275 37.885 ;
  LAYER M2 ;
        RECT 1.98 37.66 2.32 37.94 ;
  LAYER M2 ;
        RECT 6.29 37.66 6.61 37.94 ;
  LAYER M3 ;
        RECT 6.31 37.64 6.59 37.96 ;
  LAYER M2 ;
        RECT 6.29 38.08 6.61 38.36 ;
  LAYER M3 ;
        RECT 6.31 38.06 6.59 38.38 ;
  LAYER M1 ;
        RECT 2.025 37.295 2.275 37.465 ;
  LAYER M2 ;
        RECT 1.98 37.24 2.32 37.52 ;
  LAYER M1 ;
        RECT 2.025 37.715 2.275 37.885 ;
  LAYER M2 ;
        RECT 1.98 37.66 2.32 37.94 ;
  LAYER M2 ;
        RECT 6.29 37.66 6.61 37.94 ;
  LAYER M3 ;
        RECT 6.31 37.64 6.59 37.96 ;
  LAYER M2 ;
        RECT 6.29 38.08 6.61 38.36 ;
  LAYER M3 ;
        RECT 6.31 38.06 6.59 38.38 ;
  LAYER M1 ;
        RECT 2.025 37.295 2.275 37.465 ;
  LAYER M2 ;
        RECT 1.98 37.24 2.32 37.52 ;
  LAYER M1 ;
        RECT 2.025 37.715 2.275 37.885 ;
  LAYER M2 ;
        RECT 1.98 37.66 2.32 37.94 ;
  LAYER M1 ;
        RECT 8.045 37.715 8.295 37.885 ;
  LAYER M2 ;
        RECT 8 37.66 8.34 37.94 ;
  LAYER M2 ;
        RECT 6.29 37.66 6.61 37.94 ;
  LAYER M3 ;
        RECT 6.31 37.64 6.59 37.96 ;
  LAYER M2 ;
        RECT 6.29 38.08 6.61 38.36 ;
  LAYER M3 ;
        RECT 6.31 38.06 6.59 38.38 ;
  LAYER M1 ;
        RECT 2.025 37.295 2.275 37.465 ;
  LAYER M2 ;
        RECT 1.98 37.24 2.32 37.52 ;
  LAYER M1 ;
        RECT 2.025 37.715 2.275 37.885 ;
  LAYER M2 ;
        RECT 1.98 37.66 2.32 37.94 ;
  LAYER M1 ;
        RECT 8.045 37.715 8.295 37.885 ;
  LAYER M2 ;
        RECT 8 37.66 8.34 37.94 ;
  LAYER M2 ;
        RECT 6.29 37.66 6.61 37.94 ;
  LAYER M3 ;
        RECT 6.31 37.64 6.59 37.96 ;
  LAYER M2 ;
        RECT 6.29 38.08 6.61 38.36 ;
  LAYER M3 ;
        RECT 6.31 38.06 6.59 38.38 ;
  LAYER M2 ;
        RECT 1.12 33.04 2.32 33.32 ;
  LAYER M2 ;
        RECT 2.84 33.04 4.04 33.32 ;
  LAYER M2 ;
        RECT 1.12 38.08 2.32 38.36 ;
  LAYER M2 ;
        RECT 2.84 38.08 4.04 38.36 ;
  LAYER M2 ;
        RECT 6.28 34.72 7.48 35 ;
  LAYER M2 ;
        RECT 6.28 42.28 7.48 42.56 ;
  LAYER M2 ;
        RECT 2.15 33.04 3.01 33.32 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.18 2.29 38.22 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M2 ;
        RECT 2.15 38.08 3.01 38.36 ;
  LAYER M3 ;
        RECT 2.01 34.675 2.29 35.045 ;
  LAYER M2 ;
        RECT 2.15 34.72 6.45 35 ;
  LAYER M2 ;
        RECT 3.87 38.08 4.73 38.36 ;
  LAYER M1 ;
        RECT 4.605 38.22 4.855 42.42 ;
  LAYER M2 ;
        RECT 4.73 42.28 6.45 42.56 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.02 2.29 33.34 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M3 ;
        RECT 2.01 38.06 2.29 38.38 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.02 2.29 33.34 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M3 ;
        RECT 2.01 38.06 2.29 38.38 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.02 2.29 33.34 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M3 ;
        RECT 2.01 38.06 2.29 38.38 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.02 2.29 33.34 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M3 ;
        RECT 2.01 38.06 2.29 38.38 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.02 2.29 33.34 ;
  LAYER M2 ;
        RECT 1.99 34.72 2.31 35 ;
  LAYER M3 ;
        RECT 2.01 34.7 2.29 35.02 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M3 ;
        RECT 2.01 38.06 2.29 38.38 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.02 2.29 33.34 ;
  LAYER M2 ;
        RECT 1.99 34.72 2.31 35 ;
  LAYER M3 ;
        RECT 2.01 34.7 2.29 35.02 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M3 ;
        RECT 2.01 38.06 2.29 38.38 ;
  LAYER M1 ;
        RECT 4.605 38.135 4.855 38.305 ;
  LAYER M2 ;
        RECT 4.56 38.08 4.9 38.36 ;
  LAYER M1 ;
        RECT 4.605 42.335 4.855 42.505 ;
  LAYER M2 ;
        RECT 4.56 42.28 4.9 42.56 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.02 2.29 33.34 ;
  LAYER M2 ;
        RECT 1.99 34.72 2.31 35 ;
  LAYER M3 ;
        RECT 2.01 34.7 2.29 35.02 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M3 ;
        RECT 2.01 38.06 2.29 38.38 ;
  LAYER M1 ;
        RECT 4.605 38.135 4.855 38.305 ;
  LAYER M2 ;
        RECT 4.56 38.08 4.9 38.36 ;
  LAYER M1 ;
        RECT 4.605 42.335 4.855 42.505 ;
  LAYER M2 ;
        RECT 4.56 42.28 4.9 42.56 ;
  LAYER M2 ;
        RECT 1.99 33.04 2.31 33.32 ;
  LAYER M3 ;
        RECT 2.01 33.02 2.29 33.34 ;
  LAYER M2 ;
        RECT 1.99 34.72 2.31 35 ;
  LAYER M3 ;
        RECT 2.01 34.7 2.29 35.02 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M3 ;
        RECT 2.01 38.06 2.29 38.38 ;
  LAYER M1 ;
        RECT 8.905 38.135 9.155 41.665 ;
  LAYER M1 ;
        RECT 8.905 41.915 9.155 42.925 ;
  LAYER M1 ;
        RECT 8.905 44.015 9.155 45.025 ;
  LAYER M1 ;
        RECT 8.475 38.135 8.725 41.665 ;
  LAYER M1 ;
        RECT 9.335 38.135 9.585 41.665 ;
  LAYER M2 ;
        RECT 8.43 38.5 9.63 38.78 ;
  LAYER M2 ;
        RECT 8.43 44.38 9.63 44.66 ;
  LAYER M2 ;
        RECT 8 38.08 9.2 38.36 ;
  LAYER M2 ;
        RECT 8 42.28 9.2 42.56 ;
  LAYER M3 ;
        RECT 9.32 38.48 9.6 44.68 ;
  LAYER M1 ;
        RECT 8.905 33.935 9.155 37.465 ;
  LAYER M1 ;
        RECT 8.905 32.675 9.155 33.685 ;
  LAYER M1 ;
        RECT 8.905 30.575 9.155 31.585 ;
  LAYER M1 ;
        RECT 8.475 33.935 8.725 37.465 ;
  LAYER M1 ;
        RECT 9.335 33.935 9.585 37.465 ;
  LAYER M2 ;
        RECT 8.43 36.82 9.63 37.1 ;
  LAYER M2 ;
        RECT 8.43 30.94 9.63 31.22 ;
  LAYER M2 ;
        RECT 8 37.24 9.2 37.52 ;
  LAYER M2 ;
        RECT 8 33.04 9.2 33.32 ;
  LAYER M3 ;
        RECT 9.32 30.92 9.6 37.12 ;
  LAYER M1 ;
        RECT 3.745 38.135 3.995 41.665 ;
  LAYER M1 ;
        RECT 3.745 41.915 3.995 42.925 ;
  LAYER M1 ;
        RECT 3.745 44.015 3.995 45.025 ;
  LAYER M1 ;
        RECT 3.315 38.135 3.565 41.665 ;
  LAYER M1 ;
        RECT 4.175 38.135 4.425 41.665 ;
  LAYER M2 ;
        RECT 3.27 38.5 4.47 38.78 ;
  LAYER M2 ;
        RECT 3.27 44.38 4.47 44.66 ;
  LAYER M2 ;
        RECT 2.84 38.08 4.04 38.36 ;
  LAYER M2 ;
        RECT 2.84 42.28 4.04 42.56 ;
  LAYER M3 ;
        RECT 4.16 38.48 4.44 44.68 ;
  LAYER M1 ;
        RECT 6.325 38.135 6.575 41.665 ;
  LAYER M1 ;
        RECT 6.325 41.915 6.575 42.925 ;
  LAYER M1 ;
        RECT 6.325 44.015 6.575 45.025 ;
  LAYER M1 ;
        RECT 6.755 38.135 7.005 41.665 ;
  LAYER M1 ;
        RECT 5.895 38.135 6.145 41.665 ;
  LAYER M2 ;
        RECT 5.85 38.5 7.05 38.78 ;
  LAYER M2 ;
        RECT 5.85 44.38 7.05 44.66 ;
  LAYER M2 ;
        RECT 6.28 38.08 7.48 38.36 ;
  LAYER M2 ;
        RECT 6.28 42.28 7.48 42.56 ;
  LAYER M3 ;
        RECT 5.88 38.48 6.16 44.68 ;
  LAYER M1 ;
        RECT 6.325 30.575 6.575 34.105 ;
  LAYER M1 ;
        RECT 6.325 34.355 6.575 35.365 ;
  LAYER M1 ;
        RECT 6.325 36.455 6.575 37.465 ;
  LAYER M1 ;
        RECT 6.755 30.575 7.005 34.105 ;
  LAYER M1 ;
        RECT 5.895 30.575 6.145 34.105 ;
  LAYER M2 ;
        RECT 5.85 30.94 7.05 31.22 ;
  LAYER M2 ;
        RECT 5.85 36.82 7.05 37.1 ;
  LAYER M2 ;
        RECT 6.28 30.52 7.48 30.8 ;
  LAYER M2 ;
        RECT 6.28 34.72 7.48 35 ;
  LAYER M3 ;
        RECT 5.88 30.92 6.16 37.12 ;
  LAYER M1 ;
        RECT 1.165 38.135 1.415 41.665 ;
  LAYER M1 ;
        RECT 1.165 41.915 1.415 42.925 ;
  LAYER M1 ;
        RECT 1.165 44.015 1.415 45.025 ;
  LAYER M1 ;
        RECT 1.595 38.135 1.845 41.665 ;
  LAYER M1 ;
        RECT 0.735 38.135 0.985 41.665 ;
  LAYER M2 ;
        RECT 0.69 38.5 1.89 38.78 ;
  LAYER M2 ;
        RECT 0.69 44.38 1.89 44.66 ;
  LAYER M2 ;
        RECT 1.12 38.08 2.32 38.36 ;
  LAYER M2 ;
        RECT 1.12 42.28 2.32 42.56 ;
  LAYER M3 ;
        RECT 0.72 38.48 1 44.68 ;
  LAYER M1 ;
        RECT 1.165 33.935 1.415 37.465 ;
  LAYER M1 ;
        RECT 1.165 32.675 1.415 33.685 ;
  LAYER M1 ;
        RECT 1.165 30.575 1.415 31.585 ;
  LAYER M1 ;
        RECT 1.595 33.935 1.845 37.465 ;
  LAYER M1 ;
        RECT 0.735 33.935 0.985 37.465 ;
  LAYER M2 ;
        RECT 0.69 36.82 1.89 37.1 ;
  LAYER M2 ;
        RECT 0.69 30.94 1.89 31.22 ;
  LAYER M2 ;
        RECT 1.12 37.24 2.32 37.52 ;
  LAYER M2 ;
        RECT 1.12 33.04 2.32 33.32 ;
  LAYER M3 ;
        RECT 0.72 30.92 1 37.12 ;
  LAYER M1 ;
        RECT 3.745 33.935 3.995 37.465 ;
  LAYER M1 ;
        RECT 3.745 32.675 3.995 33.685 ;
  LAYER M1 ;
        RECT 3.745 30.575 3.995 31.585 ;
  LAYER M1 ;
        RECT 3.315 33.935 3.565 37.465 ;
  LAYER M1 ;
        RECT 4.175 33.935 4.425 37.465 ;
  LAYER M2 ;
        RECT 3.27 36.82 4.47 37.1 ;
  LAYER M2 ;
        RECT 3.27 30.94 4.47 31.22 ;
  LAYER M2 ;
        RECT 2.84 37.24 4.04 37.52 ;
  LAYER M2 ;
        RECT 2.84 33.04 4.04 33.32 ;
  LAYER M3 ;
        RECT 4.16 30.92 4.44 37.12 ;
  LAYER M2 ;
        RECT 1.12 22.12 2.32 22.4 ;
  LAYER M2 ;
        RECT 6.28 22.96 7.48 23.24 ;
  LAYER M2 ;
        RECT 8 17.92 9.2 18.2 ;
  LAYER M2 ;
        RECT 8 27.16 9.2 27.44 ;
  LAYER M2 ;
        RECT 8.01 17.92 8.33 18.2 ;
  LAYER M1 ;
        RECT 8.045 18.06 8.295 27.3 ;
  LAYER M2 ;
        RECT 8.01 27.16 8.33 27.44 ;
  LAYER M2 ;
        RECT 1.99 22.12 2.31 22.4 ;
  LAYER M1 ;
        RECT 2.025 22.26 2.275 22.68 ;
  LAYER M2 ;
        RECT 2.15 22.54 6.45 22.82 ;
  LAYER M3 ;
        RECT 6.31 22.68 6.59 23.1 ;
  LAYER M2 ;
        RECT 6.29 22.96 6.61 23.24 ;
  LAYER M2 ;
        RECT 6.45 22.54 8.17 22.82 ;
  LAYER M1 ;
        RECT 8.045 22.595 8.295 22.765 ;
  LAYER M1 ;
        RECT 2.025 22.175 2.275 22.345 ;
  LAYER M2 ;
        RECT 1.98 22.12 2.32 22.4 ;
  LAYER M1 ;
        RECT 2.025 22.595 2.275 22.765 ;
  LAYER M2 ;
        RECT 1.98 22.54 2.32 22.82 ;
  LAYER M2 ;
        RECT 6.29 22.54 6.61 22.82 ;
  LAYER M3 ;
        RECT 6.31 22.52 6.59 22.84 ;
  LAYER M2 ;
        RECT 6.29 22.96 6.61 23.24 ;
  LAYER M3 ;
        RECT 6.31 22.94 6.59 23.26 ;
  LAYER M1 ;
        RECT 2.025 22.175 2.275 22.345 ;
  LAYER M2 ;
        RECT 1.98 22.12 2.32 22.4 ;
  LAYER M1 ;
        RECT 2.025 22.595 2.275 22.765 ;
  LAYER M2 ;
        RECT 1.98 22.54 2.32 22.82 ;
  LAYER M2 ;
        RECT 6.29 22.54 6.61 22.82 ;
  LAYER M3 ;
        RECT 6.31 22.52 6.59 22.84 ;
  LAYER M2 ;
        RECT 6.29 22.96 6.61 23.24 ;
  LAYER M3 ;
        RECT 6.31 22.94 6.59 23.26 ;
  LAYER M1 ;
        RECT 2.025 22.175 2.275 22.345 ;
  LAYER M2 ;
        RECT 1.98 22.12 2.32 22.4 ;
  LAYER M1 ;
        RECT 2.025 22.595 2.275 22.765 ;
  LAYER M2 ;
        RECT 1.98 22.54 2.32 22.82 ;
  LAYER M1 ;
        RECT 8.045 22.595 8.295 22.765 ;
  LAYER M2 ;
        RECT 8 22.54 8.34 22.82 ;
  LAYER M2 ;
        RECT 6.29 22.54 6.61 22.82 ;
  LAYER M3 ;
        RECT 6.31 22.52 6.59 22.84 ;
  LAYER M2 ;
        RECT 6.29 22.96 6.61 23.24 ;
  LAYER M3 ;
        RECT 6.31 22.94 6.59 23.26 ;
  LAYER M1 ;
        RECT 2.025 22.175 2.275 22.345 ;
  LAYER M2 ;
        RECT 1.98 22.12 2.32 22.4 ;
  LAYER M1 ;
        RECT 2.025 22.595 2.275 22.765 ;
  LAYER M2 ;
        RECT 1.98 22.54 2.32 22.82 ;
  LAYER M1 ;
        RECT 8.045 22.595 8.295 22.765 ;
  LAYER M2 ;
        RECT 8 22.54 8.34 22.82 ;
  LAYER M2 ;
        RECT 6.29 22.54 6.61 22.82 ;
  LAYER M3 ;
        RECT 6.31 22.52 6.59 22.84 ;
  LAYER M2 ;
        RECT 6.29 22.96 6.61 23.24 ;
  LAYER M3 ;
        RECT 6.31 22.94 6.59 23.26 ;
  LAYER M2 ;
        RECT 1.12 17.92 2.32 18.2 ;
  LAYER M2 ;
        RECT 2.84 17.92 4.04 18.2 ;
  LAYER M2 ;
        RECT 1.12 22.96 2.32 23.24 ;
  LAYER M2 ;
        RECT 2.84 22.96 4.04 23.24 ;
  LAYER M2 ;
        RECT 6.28 19.6 7.48 19.88 ;
  LAYER M2 ;
        RECT 6.28 27.16 7.48 27.44 ;
  LAYER M2 ;
        RECT 2.15 17.92 3.01 18.2 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 18.06 2.29 23.1 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M2 ;
        RECT 2.15 22.96 3.01 23.24 ;
  LAYER M3 ;
        RECT 2.01 19.555 2.29 19.925 ;
  LAYER M2 ;
        RECT 2.15 19.6 6.45 19.88 ;
  LAYER M2 ;
        RECT 3.87 22.96 4.73 23.24 ;
  LAYER M1 ;
        RECT 4.605 23.1 4.855 27.3 ;
  LAYER M2 ;
        RECT 4.73 27.16 6.45 27.44 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 17.9 2.29 18.22 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.94 2.29 23.26 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 17.9 2.29 18.22 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.94 2.29 23.26 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 17.9 2.29 18.22 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.94 2.29 23.26 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 17.9 2.29 18.22 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.94 2.29 23.26 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 17.9 2.29 18.22 ;
  LAYER M2 ;
        RECT 1.99 19.6 2.31 19.88 ;
  LAYER M3 ;
        RECT 2.01 19.58 2.29 19.9 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.94 2.29 23.26 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 17.9 2.29 18.22 ;
  LAYER M2 ;
        RECT 1.99 19.6 2.31 19.88 ;
  LAYER M3 ;
        RECT 2.01 19.58 2.29 19.9 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.94 2.29 23.26 ;
  LAYER M1 ;
        RECT 4.605 23.015 4.855 23.185 ;
  LAYER M2 ;
        RECT 4.56 22.96 4.9 23.24 ;
  LAYER M1 ;
        RECT 4.605 27.215 4.855 27.385 ;
  LAYER M2 ;
        RECT 4.56 27.16 4.9 27.44 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 17.9 2.29 18.22 ;
  LAYER M2 ;
        RECT 1.99 19.6 2.31 19.88 ;
  LAYER M3 ;
        RECT 2.01 19.58 2.29 19.9 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.94 2.29 23.26 ;
  LAYER M1 ;
        RECT 4.605 23.015 4.855 23.185 ;
  LAYER M2 ;
        RECT 4.56 22.96 4.9 23.24 ;
  LAYER M1 ;
        RECT 4.605 27.215 4.855 27.385 ;
  LAYER M2 ;
        RECT 4.56 27.16 4.9 27.44 ;
  LAYER M2 ;
        RECT 1.99 17.92 2.31 18.2 ;
  LAYER M3 ;
        RECT 2.01 17.9 2.29 18.22 ;
  LAYER M2 ;
        RECT 1.99 19.6 2.31 19.88 ;
  LAYER M3 ;
        RECT 2.01 19.58 2.29 19.9 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M3 ;
        RECT 2.01 22.94 2.29 23.26 ;
  LAYER M1 ;
        RECT 8.905 23.015 9.155 26.545 ;
  LAYER M1 ;
        RECT 8.905 26.795 9.155 27.805 ;
  LAYER M1 ;
        RECT 8.905 28.895 9.155 29.905 ;
  LAYER M1 ;
        RECT 8.475 23.015 8.725 26.545 ;
  LAYER M1 ;
        RECT 9.335 23.015 9.585 26.545 ;
  LAYER M2 ;
        RECT 8.43 23.38 9.63 23.66 ;
  LAYER M2 ;
        RECT 8.43 29.26 9.63 29.54 ;
  LAYER M2 ;
        RECT 8 22.96 9.2 23.24 ;
  LAYER M2 ;
        RECT 8 27.16 9.2 27.44 ;
  LAYER M3 ;
        RECT 9.32 23.36 9.6 29.56 ;
  LAYER M1 ;
        RECT 8.905 18.815 9.155 22.345 ;
  LAYER M1 ;
        RECT 8.905 17.555 9.155 18.565 ;
  LAYER M1 ;
        RECT 8.905 15.455 9.155 16.465 ;
  LAYER M1 ;
        RECT 8.475 18.815 8.725 22.345 ;
  LAYER M1 ;
        RECT 9.335 18.815 9.585 22.345 ;
  LAYER M2 ;
        RECT 8.43 21.7 9.63 21.98 ;
  LAYER M2 ;
        RECT 8.43 15.82 9.63 16.1 ;
  LAYER M2 ;
        RECT 8 22.12 9.2 22.4 ;
  LAYER M2 ;
        RECT 8 17.92 9.2 18.2 ;
  LAYER M3 ;
        RECT 9.32 15.8 9.6 22 ;
  LAYER M1 ;
        RECT 3.745 23.015 3.995 26.545 ;
  LAYER M1 ;
        RECT 3.745 26.795 3.995 27.805 ;
  LAYER M1 ;
        RECT 3.745 28.895 3.995 29.905 ;
  LAYER M1 ;
        RECT 3.315 23.015 3.565 26.545 ;
  LAYER M1 ;
        RECT 4.175 23.015 4.425 26.545 ;
  LAYER M2 ;
        RECT 3.27 23.38 4.47 23.66 ;
  LAYER M2 ;
        RECT 3.27 29.26 4.47 29.54 ;
  LAYER M2 ;
        RECT 2.84 22.96 4.04 23.24 ;
  LAYER M2 ;
        RECT 2.84 27.16 4.04 27.44 ;
  LAYER M3 ;
        RECT 4.16 23.36 4.44 29.56 ;
  LAYER M1 ;
        RECT 6.325 23.015 6.575 26.545 ;
  LAYER M1 ;
        RECT 6.325 26.795 6.575 27.805 ;
  LAYER M1 ;
        RECT 6.325 28.895 6.575 29.905 ;
  LAYER M1 ;
        RECT 6.755 23.015 7.005 26.545 ;
  LAYER M1 ;
        RECT 5.895 23.015 6.145 26.545 ;
  LAYER M2 ;
        RECT 5.85 23.38 7.05 23.66 ;
  LAYER M2 ;
        RECT 5.85 29.26 7.05 29.54 ;
  LAYER M2 ;
        RECT 6.28 22.96 7.48 23.24 ;
  LAYER M2 ;
        RECT 6.28 27.16 7.48 27.44 ;
  LAYER M3 ;
        RECT 5.88 23.36 6.16 29.56 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 18.985 ;
  LAYER M1 ;
        RECT 6.325 19.235 6.575 20.245 ;
  LAYER M1 ;
        RECT 6.325 21.335 6.575 22.345 ;
  LAYER M1 ;
        RECT 6.755 15.455 7.005 18.985 ;
  LAYER M1 ;
        RECT 5.895 15.455 6.145 18.985 ;
  LAYER M2 ;
        RECT 5.85 15.82 7.05 16.1 ;
  LAYER M2 ;
        RECT 5.85 21.7 7.05 21.98 ;
  LAYER M2 ;
        RECT 6.28 15.4 7.48 15.68 ;
  LAYER M2 ;
        RECT 6.28 19.6 7.48 19.88 ;
  LAYER M3 ;
        RECT 5.88 15.8 6.16 22 ;
  LAYER M1 ;
        RECT 1.165 23.015 1.415 26.545 ;
  LAYER M1 ;
        RECT 1.165 26.795 1.415 27.805 ;
  LAYER M1 ;
        RECT 1.165 28.895 1.415 29.905 ;
  LAYER M1 ;
        RECT 1.595 23.015 1.845 26.545 ;
  LAYER M1 ;
        RECT 0.735 23.015 0.985 26.545 ;
  LAYER M2 ;
        RECT 0.69 23.38 1.89 23.66 ;
  LAYER M2 ;
        RECT 0.69 29.26 1.89 29.54 ;
  LAYER M2 ;
        RECT 1.12 22.96 2.32 23.24 ;
  LAYER M2 ;
        RECT 1.12 27.16 2.32 27.44 ;
  LAYER M3 ;
        RECT 0.72 23.36 1 29.56 ;
  LAYER M1 ;
        RECT 1.165 18.815 1.415 22.345 ;
  LAYER M1 ;
        RECT 1.165 17.555 1.415 18.565 ;
  LAYER M1 ;
        RECT 1.165 15.455 1.415 16.465 ;
  LAYER M1 ;
        RECT 1.595 18.815 1.845 22.345 ;
  LAYER M1 ;
        RECT 0.735 18.815 0.985 22.345 ;
  LAYER M2 ;
        RECT 0.69 21.7 1.89 21.98 ;
  LAYER M2 ;
        RECT 0.69 15.82 1.89 16.1 ;
  LAYER M2 ;
        RECT 1.12 22.12 2.32 22.4 ;
  LAYER M2 ;
        RECT 1.12 17.92 2.32 18.2 ;
  LAYER M3 ;
        RECT 0.72 15.8 1 22 ;
  LAYER M1 ;
        RECT 3.745 18.815 3.995 22.345 ;
  LAYER M1 ;
        RECT 3.745 17.555 3.995 18.565 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 16.465 ;
  LAYER M1 ;
        RECT 3.315 18.815 3.565 22.345 ;
  LAYER M1 ;
        RECT 4.175 18.815 4.425 22.345 ;
  LAYER M2 ;
        RECT 3.27 21.7 4.47 21.98 ;
  LAYER M2 ;
        RECT 3.27 15.82 4.47 16.1 ;
  LAYER M2 ;
        RECT 2.84 22.12 4.04 22.4 ;
  LAYER M2 ;
        RECT 2.84 17.92 4.04 18.2 ;
  LAYER M3 ;
        RECT 4.16 15.8 4.44 22 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M2 ;
        RECT 8.01 2.8 8.33 3.08 ;
  LAYER M1 ;
        RECT 8.045 2.94 8.295 12.18 ;
  LAYER M2 ;
        RECT 8.01 12.04 8.33 12.32 ;
  LAYER M2 ;
        RECT 1.99 7.84 2.31 8.12 ;
  LAYER M1 ;
        RECT 2.025 7.56 2.275 7.98 ;
  LAYER M2 ;
        RECT 2.15 7.42 6.45 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.14 6.59 7.56 ;
  LAYER M2 ;
        RECT 6.29 7 6.61 7.28 ;
  LAYER M2 ;
        RECT 6.45 7.42 8.17 7.7 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M1 ;
        RECT 2.025 7.475 2.275 7.645 ;
  LAYER M2 ;
        RECT 1.98 7.42 2.32 7.7 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 6.29 7 6.61 7.28 ;
  LAYER M3 ;
        RECT 6.31 6.98 6.59 7.3 ;
  LAYER M2 ;
        RECT 6.29 7.42 6.61 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.4 6.59 7.72 ;
  LAYER M1 ;
        RECT 2.025 7.475 2.275 7.645 ;
  LAYER M2 ;
        RECT 1.98 7.42 2.32 7.7 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 6.29 7 6.61 7.28 ;
  LAYER M3 ;
        RECT 6.31 6.98 6.59 7.3 ;
  LAYER M2 ;
        RECT 6.29 7.42 6.61 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.4 6.59 7.72 ;
  LAYER M1 ;
        RECT 2.025 7.475 2.275 7.645 ;
  LAYER M2 ;
        RECT 1.98 7.42 2.32 7.7 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M2 ;
        RECT 8 7.42 8.34 7.7 ;
  LAYER M2 ;
        RECT 6.29 7 6.61 7.28 ;
  LAYER M3 ;
        RECT 6.31 6.98 6.59 7.3 ;
  LAYER M2 ;
        RECT 6.29 7.42 6.61 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.4 6.59 7.72 ;
  LAYER M1 ;
        RECT 2.025 7.475 2.275 7.645 ;
  LAYER M2 ;
        RECT 1.98 7.42 2.32 7.7 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 8.045 7.475 8.295 7.645 ;
  LAYER M2 ;
        RECT 8 7.42 8.34 7.7 ;
  LAYER M2 ;
        RECT 6.29 7 6.61 7.28 ;
  LAYER M3 ;
        RECT 6.31 6.98 6.59 7.3 ;
  LAYER M2 ;
        RECT 6.29 7.42 6.61 7.7 ;
  LAYER M3 ;
        RECT 6.31 7.4 6.59 7.72 ;
  LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
  LAYER M2 ;
        RECT 2.84 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 2.15 7 3.01 7.28 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 7.14 2.29 12.18 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M2 ;
        RECT 2.15 12.04 3.01 12.32 ;
  LAYER M3 ;
        RECT 2.01 10.315 2.29 10.685 ;
  LAYER M2 ;
        RECT 2.15 10.36 6.45 10.64 ;
  LAYER M2 ;
        RECT 3.87 7 4.73 7.28 ;
  LAYER M1 ;
        RECT 4.605 2.94 4.855 7.14 ;
  LAYER M2 ;
        RECT 4.73 2.8 6.45 3.08 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 6.98 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 6.98 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 6.98 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 6.98 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 6.98 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 6.98 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M1 ;
        RECT 4.605 2.855 4.855 3.025 ;
  LAYER M2 ;
        RECT 4.56 2.8 4.9 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 6.98 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M1 ;
        RECT 4.605 2.855 4.855 3.025 ;
  LAYER M2 ;
        RECT 4.56 2.8 4.9 3.08 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
  LAYER M3 ;
        RECT 2.01 6.98 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.99 10.36 2.31 10.64 ;
  LAYER M3 ;
        RECT 2.01 10.34 2.29 10.66 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M3 ;
        RECT 2.01 12.02 2.29 12.34 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 8 7 9.2 7.28 ;
  LAYER M2 ;
        RECT 8 2.8 9.2 3.08 ;
  LAYER M3 ;
        RECT 9.32 0.68 9.6 6.88 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 8.43 14.14 9.63 14.42 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 2.84 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 2.84 2.8 4.04 3.08 ;
  LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M2 ;
        RECT 5.85 6.58 7.05 6.86 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 6.88 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M3 ;
        RECT 0.72 0.68 1 6.88 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M3 ;
        RECT 0.72 8.24 1 14.44 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  LAYER M4 ;
        RECT 11.18 1.67 18.48 8.97 ;
  LAYER M4 ;
        RECT 18.03 1.46 18.48 3.98 ;
  LAYER M5 ;
        RECT 11.405 7.99 11.855 10.51 ;
  LAYER M4 ;
        RECT 10.585 9.68 18.225 10.48 ;
  LAYER M4 ;
        RECT 10.585 0.86 18.225 1.66 ;
  LAYER M4 ;
        RECT 11.18 13.01 18.48 20.31 ;
  LAYER M4 ;
        RECT 18.03 12.8 18.48 15.32 ;
  LAYER M5 ;
        RECT 11.405 19.33 11.855 21.85 ;
  LAYER M4 ;
        RECT 10.585 21.02 18.225 21.82 ;
  LAYER M4 ;
        RECT 10.585 12.2 18.225 13 ;
  LAYER M4 ;
        RECT 11.18 24.35 18.48 31.65 ;
  LAYER M4 ;
        RECT 18.03 24.14 18.48 26.66 ;
  LAYER M5 ;
        RECT 11.405 30.67 11.855 33.19 ;
  LAYER M4 ;
        RECT 10.585 32.36 18.225 33.16 ;
  LAYER M4 ;
        RECT 10.585 23.54 18.225 24.34 ;
  LAYER M4 ;
        RECT 11.18 35.69 18.48 42.99 ;
  LAYER M4 ;
        RECT 18.03 35.48 18.48 38 ;
  LAYER M5 ;
        RECT 11.405 42.01 11.855 44.53 ;
  LAYER M4 ;
        RECT 10.585 43.7 18.225 44.5 ;
  LAYER M4 ;
        RECT 10.585 34.88 18.225 35.68 ;
  END 
END TWO_BIT_RES_DAC
