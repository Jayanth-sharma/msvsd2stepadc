magic
tech sky130A
magscale 1 2
timestamp 1679679491
<< locali >>
rect 405 2419 413 2453
rect 447 2419 455 2453
rect 405 2369 455 2419
rect 405 2335 413 2369
rect 447 2335 455 2369
rect 577 2335 585 2369
rect 619 2335 627 2369
rect 577 1613 627 2335
rect 577 1579 585 1613
rect 619 1579 627 1613
rect 577 1445 627 1579
rect 577 1411 585 1445
rect 619 1411 627 1445
rect 577 1277 627 1411
rect 405 1243 413 1277
rect 447 1243 455 1277
rect 577 1243 585 1277
rect 619 1243 627 1277
rect 405 605 455 1243
rect 405 571 413 605
rect 447 571 455 605
<< viali >>
rect 413 2419 447 2453
rect 413 2335 447 2369
rect 585 2335 619 2369
rect 585 1579 619 1613
rect 585 1411 619 1445
rect 413 1243 447 1277
rect 585 1243 619 1277
rect 413 571 447 605
<< metal1 >>
rect 396 2453 464 2464
rect 396 2419 413 2453
rect 447 2419 464 2453
rect 396 2408 464 2419
rect 656 2462 720 2464
rect 656 2410 662 2462
rect 714 2410 720 2462
rect 656 2408 720 2410
rect 396 2369 636 2380
rect 396 2335 413 2369
rect 447 2335 585 2369
rect 619 2335 636 2369
rect 396 2324 636 2335
rect 312 1622 376 1624
rect 312 1570 318 1622
rect 370 1570 376 1622
rect 312 1568 376 1570
rect 568 1613 636 1624
rect 568 1579 585 1613
rect 619 1579 636 1613
rect 568 1568 636 1579
rect 312 1454 376 1456
rect 312 1402 318 1454
rect 370 1402 376 1454
rect 312 1400 376 1402
rect 568 1445 636 1456
rect 568 1411 585 1445
rect 619 1411 636 1445
rect 568 1400 636 1411
rect 396 1277 636 1288
rect 396 1243 413 1277
rect 447 1243 585 1277
rect 619 1243 636 1277
rect 396 1232 636 1243
rect 396 605 464 616
rect 396 571 413 605
rect 447 571 464 605
rect 396 560 464 571
rect 656 614 720 616
rect 656 562 662 614
rect 714 562 720 614
rect 656 560 720 562
<< via1 >>
rect 662 2410 714 2462
rect 318 1570 370 1622
rect 318 1402 370 1454
rect 662 562 714 614
<< metal2 >>
rect 660 2462 716 2468
rect 660 2410 662 2462
rect 714 2410 716 2462
rect 316 1622 372 1628
rect 316 1570 318 1622
rect 370 1570 372 1622
rect 316 1454 372 1570
rect 316 1402 318 1454
rect 370 1402 372 1454
rect 316 1396 372 1402
rect 660 614 716 2410
rect 660 562 662 614
rect 714 562 716 614
rect 660 556 716 562
use NMOS_S_42092372_X1_Y1_1679678942_1679678944  NMOS_S_42092372_X1_Y1_1679678942_1679678944_0
timestamp 1679679491
transform -1 0 516 0 -1 1512
box 52 56 395 1482
use NMOS_S_42092372_X1_Y1_1679678942_1679678944  NMOS_S_42092372_X1_Y1_1679678942_1679678944_1
timestamp 1679679491
transform 1 0 516 0 -1 1512
box 52 56 395 1482
use PMOS_S_45039047_X1_Y1_1679678943_1679678944  PMOS_S_45039047_X1_Y1_1679678943_1679678944_0
timestamp 1679679491
transform -1 0 516 0 1 1512
box 0 0 516 1512
use PMOS_S_45039047_X1_Y1_1679678943_1679678944  PMOS_S_45039047_X1_Y1_1679678943_1679678944_1
timestamp 1679679491
transform 1 0 516 0 1 1512
box 0 0 516 1512
<< end >>
