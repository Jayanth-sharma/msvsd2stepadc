* SPICE3 file created from RING_OSC_0.ext - technology: sky130A
.option scale=5000u
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
V1 VDD GND 1.8

x1 VDD Y GND ring_osc

**** begin user architecture code



* .dc V2 0 1.8 0.01
.tran 10p 4n 0
.control
  run
  print allv > plot_data_v.txt
  print alli > plot_data_i.txt
  plot v(Y)
.endc



**** end user architecture code

.subckt ring_osc VDD Y GND
X0 m1_688_4424# li_405_1579# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=6.678e+11p ps=8.22e+06u w=420000u l=150000u
X1 VSUBS li_405_1579# m1_688_4424# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 m1_688_4424# li_405_1579# m1_398_2912# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=6.678e+11p ps=8.22e+06u w=420000u l=150000u
X3 m1_398_2912# li_405_1579# m1_688_4424# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 li_405_1579# STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# m1_398_2912# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X5 m1_398_2912# STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# li_405_1579# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# m1_688_4424# m1_398_2912# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X7 m1_398_2912# m1_688_4424# STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 li_405_1579# STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X9 VSUBS STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# li_405_1579# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# m1_688_4424# VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X11 Y m1_688_4424# STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 m1_688_4424# m1_398_2912# 2.28fF
C1 Y li_405_1579# 0.01fF
C2 GND Y 0.02fF
C3 VDD STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# 0.03fF
C4 li_405_1579# STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# 0.59fF
C5 m1_398_2912# STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# 2.97fF
C6 li_405_1579# VDD 1.31fF
C7 GND STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# 0.15fF
C8 m1_688_4424# STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# 0.62fF
C9 GND VDD 0.24fF
C10 m1_688_4424# VDD 0.32fF
C11 Y STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# 0.00fF
C12 li_405_1579# m1_398_2912# 2.12fF
C13 Y VDD 0.24fF
C14 GND li_405_1579# 0.14fF
C15 m1_688_4424# li_405_1579# 0.46fF
C16 VDD VSUBS 0.16fF
C17 m1_688_4424# VSUBS 2.58fF
C18 li_405_1579# VSUBS 1.88fF 
C19 STAGE2_INV_5734008_0_0_1677844589_0/li_491_571# VSUBS 1.16fF 
C20 m1_398_2912# VSUBS 8.15fF
.ends


