magic
tech sky130A
magscale 1 2
timestamp 1678186317
<< locali >>
rect 128 500 1182 508
rect 172 498 1182 500
rect 172 442 1126 498
rect 1174 442 1182 498
<< viali >>
rect 128 442 172 500
rect 1126 440 1174 498
<< metal1 >>
rect -52 1108 1202 1274
rect -20 956 24 1108
rect 128 1002 192 1062
rect -20 862 134 956
rect 388 950 430 1108
rect 536 1000 598 1056
rect 810 960 848 1108
rect 952 1010 1014 1066
rect 182 778 336 880
rect 388 848 540 950
rect 128 720 190 730
rect 122 674 190 720
rect 122 500 178 674
rect 122 442 128 500
rect 172 442 178 500
rect 122 284 178 442
rect 288 496 332 778
rect 596 772 746 898
rect 810 848 958 960
rect 1106 910 1162 912
rect 1012 784 1162 910
rect 536 672 598 728
rect 544 496 594 672
rect 288 452 594 496
rect 118 228 180 284
rect 288 186 332 452
rect 544 278 594 452
rect 712 498 746 772
rect 968 738 1014 744
rect 952 682 1014 738
rect 968 498 1014 682
rect 712 454 1014 498
rect 544 224 606 278
rect 712 188 746 454
rect 968 274 1014 454
rect 1106 518 1162 784
rect 1106 498 1258 518
rect 1106 440 1126 498
rect 1174 440 1258 498
rect 1106 434 1258 440
rect 964 220 1026 274
rect -24 98 12 102
rect -30 4 122 98
rect 172 80 332 186
rect 288 78 332 80
rect 400 4 552 98
rect 598 64 756 188
rect 1106 180 1162 434
rect 820 98 856 102
rect 712 60 746 64
rect 818 4 970 98
rect 1018 54 1168 180
rect 1106 52 1162 54
rect -24 -140 12 4
rect 116 -82 180 -30
rect 402 -140 438 4
rect 544 -90 606 -34
rect 820 -140 856 4
rect 964 -92 1026 -38
rect -60 -280 1188 -140
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1678186317
transform 1 0 158 0 1 866
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1678186317
transform 1 0 567 0 1 865
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 1678186317
transform 1 0 983 0 1 873
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1678186317
transform 1 0 575 0 1 94
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 1678186317
transform 1 0 148 0 1 99
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM6
timestamp 1678186317
transform 1 0 995 0 1 90
box -211 -310 211 310
<< labels >>
rlabel metal1 1134 1114 1200 1272 3 vp
port 1 e
rlabel metal1 1184 434 1258 518 3 y
port 2 e
rlabel metal1 1114 -280 1188 -196 3 vn
port 3 e
<< end >>
