magic
tech sky130A
magscale 1 2
timestamp 1679679491
<< nwell >>
rect 0 0 516 1512
<< pmos >>
rect 200 315 230 819
rect 286 315 316 819
<< pdiff >>
rect 147 705 200 819
rect 147 671 155 705
rect 189 671 200 705
rect 147 637 200 671
rect 147 603 155 637
rect 189 603 200 637
rect 147 569 200 603
rect 147 535 155 569
rect 189 535 200 569
rect 147 501 200 535
rect 147 467 155 501
rect 189 467 200 501
rect 147 433 200 467
rect 147 399 155 433
rect 189 399 200 433
rect 147 365 200 399
rect 147 331 155 365
rect 189 331 200 365
rect 147 315 200 331
rect 230 705 286 819
rect 230 671 241 705
rect 275 671 286 705
rect 230 637 286 671
rect 230 603 241 637
rect 275 603 286 637
rect 230 569 286 603
rect 230 535 241 569
rect 275 535 286 569
rect 230 501 286 535
rect 230 467 241 501
rect 275 467 286 501
rect 230 433 286 467
rect 230 399 241 433
rect 275 399 286 433
rect 230 365 286 399
rect 230 331 241 365
rect 275 331 286 365
rect 230 315 286 331
rect 316 705 369 819
rect 316 671 327 705
rect 361 671 369 705
rect 316 637 369 671
rect 316 603 327 637
rect 361 603 369 637
rect 316 569 369 603
rect 316 535 327 569
rect 361 535 369 569
rect 316 501 369 535
rect 316 467 327 501
rect 361 467 369 501
rect 316 433 369 467
rect 316 399 327 433
rect 361 399 369 433
rect 316 365 369 399
rect 316 331 327 365
rect 361 331 369 365
rect 316 315 369 331
<< pdiffc >>
rect 155 671 189 705
rect 155 603 189 637
rect 155 535 189 569
rect 155 467 189 501
rect 155 399 189 433
rect 155 331 189 365
rect 241 671 275 705
rect 241 603 275 637
rect 241 535 275 569
rect 241 467 275 501
rect 241 399 275 433
rect 241 331 275 365
rect 327 671 361 705
rect 327 603 361 637
rect 327 535 361 569
rect 327 467 361 501
rect 327 399 361 433
rect 327 331 361 365
<< nsubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
<< nsubdiffcont >>
rect 241 1327 275 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 819 230 897
rect 286 819 316 897
rect 200 252 230 315
rect 286 252 316 315
<< polycont >>
rect 241 907 275 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 147 705 197 773
rect 147 671 155 705
rect 189 671 197 705
rect 147 637 197 671
rect 147 603 155 637
rect 189 603 197 637
rect 147 569 197 603
rect 147 535 155 569
rect 189 535 197 569
rect 147 501 197 535
rect 147 467 155 501
rect 189 467 197 501
rect 147 433 197 467
rect 147 399 155 433
rect 189 399 197 433
rect 147 365 197 399
rect 147 331 155 365
rect 189 331 197 365
rect 147 185 197 331
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 705 283 773
rect 233 671 241 705
rect 275 671 283 705
rect 233 637 283 671
rect 233 603 241 637
rect 275 603 283 637
rect 233 569 283 603
rect 233 535 241 569
rect 275 535 283 569
rect 233 501 283 535
rect 233 467 241 501
rect 275 467 283 501
rect 233 433 283 467
rect 233 399 241 433
rect 275 399 283 433
rect 233 365 283 399
rect 233 331 241 365
rect 275 331 283 365
rect 233 101 283 331
rect 233 67 241 101
rect 275 67 283 101
rect 319 705 369 773
rect 319 671 327 705
rect 361 671 369 705
rect 319 637 369 671
rect 319 603 327 637
rect 361 603 369 637
rect 319 569 369 603
rect 319 535 327 569
rect 361 535 369 569
rect 319 501 369 535
rect 319 467 327 501
rect 361 467 369 501
rect 319 433 369 467
rect 319 399 327 433
rect 361 399 369 433
rect 319 365 369 399
rect 319 331 327 365
rect 361 331 369 365
rect 319 185 369 331
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
<< viali >>
rect 241 1327 275 1361
rect 241 907 275 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
<< metal1 >>
rect 138 1370 378 1372
rect 138 1361 318 1370
rect 138 1327 241 1361
rect 275 1327 318 1361
rect 138 1318 318 1327
rect 370 1318 378 1370
rect 138 1316 378 1318
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 194 378 196
rect 138 185 318 194
rect 138 151 155 185
rect 189 151 318 185
rect 138 142 318 151
rect 370 142 378 194
rect 138 140 378 142
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< via1 >>
rect 318 1318 370 1370
rect 318 185 370 194
rect 318 151 327 185
rect 327 151 361 185
rect 361 151 370 185
rect 318 142 370 151
<< metal2 >>
rect 316 1370 372 1376
rect 316 1318 318 1370
rect 370 1318 372 1370
rect 316 194 372 1318
rect 316 142 318 194
rect 370 142 372 194
rect 316 136 372 142
<< end >>
