** sch_path: /home/vinayreddy/Desktop/mspdr/week7/pre-layout/tb_2bitADC.sch
**.subckt tb_2bitADC b3 b2 b1 Vb Vref Vin VCC
*.opin b3
*.opin b2
*.opin b1
*.ipin Vb
*.ipin Vref
*.ipin Vin
*.iopin VCC
x1 Vref Vin VCC Vb b3 b2 b1 GND Two_BitADC
V1 VCC GND 3.3
.save i(v1)
V2 Vb GND 0.9
.save i(v2)
V3 Vref GND sine(0 3.3 10000000)
.save i(v3)
V4 Vin GND 4.2
.save i(v4)
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 10p 100n
.control
run
save all
.endc

**** end user architecture code
**.ends

* expanding   symbol:  Two_BitADC.sym # of pins=8
** sym_path: /home/vinayreddy/Desktop/mspdr/week7/pre-layout/Two_BitADC.sym
** sch_path: /home/vinayreddy/Desktop/mspdr/week7/pre-layout/Two_BitADC.sch
.subckt Two_BitADC INN INP VCC BIAS C3 C2 C1 GND
*.iopin VCC
*.ipin BIAS
*.opin C3
*.opin C2
*.opin C1
*.ipin INN
*.ipin INP
*.iopin GND
x1 VCC C3 net1 INN GND BIAS comp
XR1 net1 INP INP sky130_fd_pr__res_generic_pd W=10 L=5.2 mult=1 m=1
XR2 net2 net1 net1 sky130_fd_pr__res_generic_pd W=10 L=5.2 mult=1 m=1
XR3 net3 net2 net2 sky130_fd_pr__res_generic_pd W=10 L=5.2 mult=1 m=1
XR4 GND net3 net3 sky130_fd_pr__res_generic_pd W=10 L=5.2 mult=1 m=1
x2 VCC C2 net2 INN GND BIAS comp
x3 VCC C1 net3 INN GND BIAS comp
.ends


* expanding   symbol:  comp.sym # of pins=6
** sym_path: /home/vinayreddy/Desktop/mspdr/week7/pre-layout/comp.sym
** sch_path: /home/vinayreddy/Desktop/mspdr/week7/pre-layout/comp.sch
.subckt comp VCC OUT INN INP GND BIAS
*.ipin BIAS
*.iopin VCC
*.iopin GND
*.opin OUT
*.ipin INN
*.ipin INP
XM1 net3 net3 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 INN net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 net1 BIAS GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 net3 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 INP net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 net2 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net4 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 net5 net4 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 OUT net5 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 net5 net4 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 OUT net5 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
