** sch_path: /home/vinayreddy/Desktop/mspdr/ALIGN-public/work/inv_tb.sch
**.subckt inv_tb out in
*.opin out
*.ipin in
x1 net1 in out GND inv
V1 net1 GND 1.8
.save i(v1)
V2 in GND pulse(0 1.8 1n 1n 1n 2n 4n)
.save i(v2)
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 0.01n 20n
.save all


**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/vinayreddy/Desktop/mspdr/ALIGN-public/work/inv.sym
** sch_path: /home/vinayreddy/Desktop/mspdr/ALIGN-public/work/inv.sch
.subckt inv Vdd! Vin Vout Vss!
*.ipin Vin
*.opin Vout
*.iopin Vdd!
*.iopin Vss!
XM1 Vout Vin Vdd! Vdd! sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin Vss! Vss! sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
