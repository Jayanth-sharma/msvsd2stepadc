MACRO TWO_BIT_RES_DAC
  ORIGIN 0 0 ;
  FOREIGN TWO_BIT_RES_DAC 0 0 ;
  SIZE 20.8 BY 50.99 ;
  PIN D0
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 17.08 2.32 17.36 ;
      LAYER M2 ;
        RECT 2.84 17.08 4.04 17.36 ;
      LAYER M2 ;
        RECT 2.15 17.08 3.01 17.36 ;
      LAYER M2 ;
        RECT 1.12 47.32 2.32 47.6 ;
      LAYER M2 ;
        RECT 2.84 47.32 4.04 47.6 ;
      LAYER M2 ;
        RECT 2.15 47.32 3.01 47.6 ;
      LAYER M2 ;
        RECT 2.42 17.08 2.74 17.36 ;
      LAYER M3 ;
        RECT 2.44 17.22 2.72 47.46 ;
      LAYER M2 ;
        RECT 2.42 47.32 2.74 47.6 ;
    END
  END D0
  PIN INP2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 9.32 43.52 9.6 49.72 ;
      LAYER M2 ;
        RECT 6.28 49.84 7.48 50.12 ;
      LAYER M3 ;
        RECT 9.32 49.56 9.6 49.98 ;
      LAYER M2 ;
        RECT 7.31 49.84 9.46 50.12 ;
      LAYER M4 ;
        RECT 10.585 48.74 19.515 49.54 ;
      LAYER M3 ;
        RECT 9.32 48.955 9.6 49.325 ;
      LAYER M4 ;
        RECT 9.46 48.74 10.75 49.54 ;
    END
  END INP2
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 32.2 2.32 32.48 ;
      LAYER M2 ;
        RECT 2.84 32.2 4.04 32.48 ;
      LAYER M2 ;
        RECT 2.15 32.2 3.01 32.48 ;
    END
  END D1
  PIN OUT_V
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 5.88 20.84 6.16 27.04 ;
      LAYER M2 ;
        RECT 8 27.16 9.2 27.44 ;
      LAYER M2 ;
        RECT 8 28 9.2 28.28 ;
      LAYER M2 ;
        RECT 8.44 27.16 8.76 27.44 ;
      LAYER M3 ;
        RECT 8.46 27.3 8.74 28.14 ;
      LAYER M2 ;
        RECT 8.44 28 8.76 28.28 ;
      LAYER M3 ;
        RECT 5.88 28.4 6.16 34.6 ;
      LAYER M3 ;
        RECT 5.88 26.275 6.16 26.645 ;
      LAYER M4 ;
        RECT 6.02 26.06 8.17 26.86 ;
      LAYER M3 ;
        RECT 8.03 26.46 8.31 27.3 ;
      LAYER M2 ;
        RECT 8.01 27.16 8.33 27.44 ;
      LAYER M3 ;
        RECT 5.88 26.88 6.16 28.56 ;
    END
  END OUT_V
  PIN INP1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 10.585 0.86 19.515 1.66 ;
    END
  END INP1
  OBS 
  LAYER M3 ;
        RECT 9.32 35.96 9.6 42.16 ;
  LAYER M2 ;
        RECT 6.28 42.28 7.48 42.56 ;
  LAYER M3 ;
        RECT 9.32 41.395 9.6 41.765 ;
  LAYER M2 ;
        RECT 7.31 41.44 9.46 41.72 ;
  LAYER M1 ;
        RECT 7.185 41.58 7.435 42.42 ;
  LAYER M2 ;
        RECT 7.15 42.28 7.47 42.56 ;
  LAYER M4 ;
        RECT 10.585 36.14 19.515 36.94 ;
  LAYER M4 ;
        RECT 10.585 38.66 19.515 39.46 ;
  LAYER M4 ;
        RECT 14.885 36.14 15.215 36.94 ;
  LAYER M3 ;
        RECT 14.91 36.54 15.19 39.06 ;
  LAYER M4 ;
        RECT 14.885 38.66 15.215 39.46 ;
  LAYER M3 ;
        RECT 9.32 38.875 9.6 39.245 ;
  LAYER M4 ;
        RECT 9.46 38.66 10.75 39.46 ;
  LAYER M3 ;
        RECT 9.32 38.875 9.6 39.245 ;
  LAYER M4 ;
        RECT 9.295 38.66 9.625 39.46 ;
  LAYER M3 ;
        RECT 9.32 38.875 9.6 39.245 ;
  LAYER M4 ;
        RECT 9.295 38.66 9.625 39.46 ;
  LAYER M3 ;
        RECT 9.32 28.4 9.6 34.6 ;
  LAYER M2 ;
        RECT 6.28 34.72 7.48 35 ;
  LAYER M3 ;
        RECT 9.32 34.44 9.6 34.86 ;
  LAYER M2 ;
        RECT 7.31 34.72 9.46 35 ;
  LAYER M3 ;
        RECT 5.88 35.96 6.16 42.16 ;
  LAYER M2 ;
        RECT 8 42.28 9.2 42.56 ;
  LAYER M2 ;
        RECT 8 43.12 9.2 43.4 ;
  LAYER M2 ;
        RECT 8.44 42.28 8.76 42.56 ;
  LAYER M3 ;
        RECT 8.46 42.42 8.74 43.26 ;
  LAYER M2 ;
        RECT 8.44 43.12 8.76 43.4 ;
  LAYER M3 ;
        RECT 5.88 43.52 6.16 49.72 ;
  LAYER M3 ;
        RECT 5.88 41.395 6.16 41.765 ;
  LAYER M4 ;
        RECT 6.02 41.18 8.17 41.98 ;
  LAYER M3 ;
        RECT 8.03 41.58 8.31 42.42 ;
  LAYER M2 ;
        RECT 8.01 42.28 8.33 42.56 ;
  LAYER M3 ;
        RECT 5.88 42 6.16 43.68 ;
  LAYER M2 ;
        RECT 6.29 34.72 6.61 35 ;
  LAYER M3 ;
        RECT 6.31 34.86 6.59 35.7 ;
  LAYER M2 ;
        RECT 6.02 35.56 6.45 35.84 ;
  LAYER M3 ;
        RECT 5.88 35.7 6.16 36.12 ;
  LAYER M2 ;
        RECT 5.86 35.56 6.18 35.84 ;
  LAYER M3 ;
        RECT 5.88 35.54 6.16 35.86 ;
  LAYER M2 ;
        RECT 6.29 34.72 6.61 35 ;
  LAYER M3 ;
        RECT 6.31 34.7 6.59 35.02 ;
  LAYER M2 ;
        RECT 6.29 35.56 6.61 35.84 ;
  LAYER M3 ;
        RECT 6.31 35.54 6.59 35.86 ;
  LAYER M2 ;
        RECT 5.86 35.56 6.18 35.84 ;
  LAYER M3 ;
        RECT 5.88 35.54 6.16 35.86 ;
  LAYER M2 ;
        RECT 6.29 34.72 6.61 35 ;
  LAYER M3 ;
        RECT 6.31 34.7 6.59 35.02 ;
  LAYER M2 ;
        RECT 6.29 35.56 6.61 35.84 ;
  LAYER M3 ;
        RECT 6.31 35.54 6.59 35.86 ;
  LAYER M3 ;
        RECT 9.32 5.72 9.6 11.92 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M3 ;
        RECT 9.32 11.155 9.6 11.525 ;
  LAYER M2 ;
        RECT 7.31 11.2 9.46 11.48 ;
  LAYER M1 ;
        RECT 7.185 11.34 7.435 12.18 ;
  LAYER M2 ;
        RECT 7.15 12.04 7.47 12.32 ;
  LAYER M4 ;
        RECT 10.585 10.94 19.515 11.74 ;
  LAYER M4 ;
        RECT 10.585 13.46 19.515 14.26 ;
  LAYER M4 ;
        RECT 14.885 10.94 15.215 11.74 ;
  LAYER M3 ;
        RECT 14.91 11.34 15.19 13.86 ;
  LAYER M4 ;
        RECT 14.885 13.46 15.215 14.26 ;
  LAYER M2 ;
        RECT 9.46 11.2 10.75 11.48 ;
  LAYER M3 ;
        RECT 10.61 11.219 10.89 11.461 ;
  LAYER M4 ;
        RECT 10.585 10.94 10.915 11.74 ;
  LAYER M2 ;
        RECT 10.59 11.2 10.91 11.48 ;
  LAYER M3 ;
        RECT 10.61 11.18 10.89 11.5 ;
  LAYER M3 ;
        RECT 10.61 11.155 10.89 11.525 ;
  LAYER M4 ;
        RECT 10.585 10.94 10.915 11.74 ;
  LAYER M3 ;
        RECT 9.32 13.28 9.6 19.48 ;
  LAYER M2 ;
        RECT 6.28 19.6 7.48 19.88 ;
  LAYER M3 ;
        RECT 9.32 19.32 9.6 19.74 ;
  LAYER M2 ;
        RECT 7.31 19.6 9.46 19.88 ;
  LAYER M4 ;
        RECT 10.585 23.54 19.515 24.34 ;
  LAYER M4 ;
        RECT 10.585 26.06 19.515 26.86 ;
  LAYER M2 ;
        RECT 9.46 19.6 10.75 19.88 ;
  LAYER M3 ;
        RECT 10.61 19.74 10.89 23.94 ;
  LAYER M4 ;
        RECT 10.585 23.54 10.915 24.34 ;
  LAYER M3 ;
        RECT 10.61 23.94 10.89 26.46 ;
  LAYER M4 ;
        RECT 10.585 26.06 10.915 26.86 ;
  LAYER M2 ;
        RECT 10.59 19.6 10.91 19.88 ;
  LAYER M3 ;
        RECT 10.61 19.58 10.89 19.9 ;
  LAYER M3 ;
        RECT 10.61 23.755 10.89 24.125 ;
  LAYER M4 ;
        RECT 10.585 23.54 10.915 24.34 ;
  LAYER M2 ;
        RECT 10.59 19.6 10.91 19.88 ;
  LAYER M3 ;
        RECT 10.61 19.58 10.89 19.9 ;
  LAYER M3 ;
        RECT 10.61 23.755 10.89 24.125 ;
  LAYER M4 ;
        RECT 10.585 23.54 10.915 24.34 ;
  LAYER M2 ;
        RECT 10.59 19.6 10.91 19.88 ;
  LAYER M3 ;
        RECT 10.61 19.58 10.89 19.9 ;
  LAYER M3 ;
        RECT 10.61 23.755 10.89 24.125 ;
  LAYER M4 ;
        RECT 10.585 23.54 10.915 24.34 ;
  LAYER M3 ;
        RECT 10.61 26.275 10.89 26.645 ;
  LAYER M4 ;
        RECT 10.585 26.06 10.915 26.86 ;
  LAYER M2 ;
        RECT 10.59 19.6 10.91 19.88 ;
  LAYER M3 ;
        RECT 10.61 19.58 10.89 19.9 ;
  LAYER M3 ;
        RECT 10.61 23.755 10.89 24.125 ;
  LAYER M4 ;
        RECT 10.585 23.54 10.915 24.34 ;
  LAYER M3 ;
        RECT 10.61 26.275 10.89 26.645 ;
  LAYER M4 ;
        RECT 10.585 26.06 10.915 26.86 ;
  LAYER M3 ;
        RECT 5.88 5.72 6.16 11.92 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M2 ;
        RECT 8 12.88 9.2 13.16 ;
  LAYER M2 ;
        RECT 8.44 12.04 8.76 12.32 ;
  LAYER M3 ;
        RECT 8.46 12.18 8.74 13.02 ;
  LAYER M2 ;
        RECT 8.44 12.88 8.76 13.16 ;
  LAYER M3 ;
        RECT 5.88 13.28 6.16 19.48 ;
  LAYER M3 ;
        RECT 5.88 11.155 6.16 11.525 ;
  LAYER M4 ;
        RECT 6.02 10.94 8.17 11.74 ;
  LAYER M3 ;
        RECT 8.03 11.34 8.31 12.18 ;
  LAYER M2 ;
        RECT 8.01 12.04 8.33 12.32 ;
  LAYER M3 ;
        RECT 5.88 11.76 6.16 13.44 ;
  LAYER M3 ;
        RECT 9.32 20.84 9.6 27.04 ;
  LAYER M2 ;
        RECT 6.28 27.16 7.48 27.44 ;
  LAYER M3 ;
        RECT 9.32 26.275 9.6 26.645 ;
  LAYER M2 ;
        RECT 7.31 26.32 9.46 26.6 ;
  LAYER M1 ;
        RECT 7.185 26.46 7.435 27.3 ;
  LAYER M2 ;
        RECT 7.15 27.16 7.47 27.44 ;
  LAYER M3 ;
        RECT 5.88 19.32 6.16 20.16 ;
  LAYER M2 ;
        RECT 6.02 20.02 9.46 20.3 ;
  LAYER M1 ;
        RECT 9.335 20.16 9.585 20.58 ;
  LAYER M2 ;
        RECT 9.311 20.44 9.609 20.72 ;
  LAYER M3 ;
        RECT 9.32 20.58 9.6 21 ;
  LAYER M1 ;
        RECT 9.335 20.075 9.585 20.245 ;
  LAYER M2 ;
        RECT 9.29 20.02 9.63 20.3 ;
  LAYER M1 ;
        RECT 9.335 20.495 9.585 20.665 ;
  LAYER M2 ;
        RECT 9.29 20.44 9.63 20.72 ;
  LAYER M2 ;
        RECT 5.86 20.02 6.18 20.3 ;
  LAYER M3 ;
        RECT 5.88 20 6.16 20.32 ;
  LAYER M2 ;
        RECT 9.3 20.44 9.62 20.72 ;
  LAYER M3 ;
        RECT 9.32 20.42 9.6 20.74 ;
  LAYER M1 ;
        RECT 9.335 20.075 9.585 20.245 ;
  LAYER M2 ;
        RECT 9.29 20.02 9.63 20.3 ;
  LAYER M2 ;
        RECT 5.86 20.02 6.18 20.3 ;
  LAYER M3 ;
        RECT 5.88 20 6.16 20.32 ;
  LAYER M2 ;
        RECT 1.12 42.28 2.32 42.56 ;
  LAYER M2 ;
        RECT 3.7 42.28 4.9 42.56 ;
  LAYER M2 ;
        RECT 8 38.08 9.2 38.36 ;
  LAYER M2 ;
        RECT 8 47.32 9.2 47.6 ;
  LAYER M2 ;
        RECT 8.01 38.08 8.33 38.36 ;
  LAYER M1 ;
        RECT 8.045 38.22 8.295 47.46 ;
  LAYER M2 ;
        RECT 8.01 47.32 8.33 47.6 ;
  LAYER M2 ;
        RECT 2.15 42.28 3.87 42.56 ;
  LAYER M2 ;
        RECT 4.73 42.28 5.59 42.56 ;
  LAYER M1 ;
        RECT 5.465 42.42 5.715 42.84 ;
  LAYER M2 ;
        RECT 5.59 42.7 8.17 42.98 ;
  LAYER M1 ;
        RECT 8.045 42.755 8.295 42.925 ;
  LAYER M1 ;
        RECT 5.465 42.335 5.715 42.505 ;
  LAYER M2 ;
        RECT 5.42 42.28 5.76 42.56 ;
  LAYER M1 ;
        RECT 5.465 42.755 5.715 42.925 ;
  LAYER M2 ;
        RECT 5.42 42.7 5.76 42.98 ;
  LAYER M1 ;
        RECT 8.045 42.755 8.295 42.925 ;
  LAYER M2 ;
        RECT 8 42.7 8.34 42.98 ;
  LAYER M1 ;
        RECT 5.465 42.335 5.715 42.505 ;
  LAYER M2 ;
        RECT 5.42 42.28 5.76 42.56 ;
  LAYER M1 ;
        RECT 5.465 42.755 5.715 42.925 ;
  LAYER M2 ;
        RECT 5.42 42.7 5.76 42.98 ;
  LAYER M1 ;
        RECT 8.045 42.755 8.295 42.925 ;
  LAYER M2 ;
        RECT 8 42.7 8.34 42.98 ;
  LAYER M2 ;
        RECT 1.12 38.08 2.32 38.36 ;
  LAYER M2 ;
        RECT 3.7 38.08 4.9 38.36 ;
  LAYER M2 ;
        RECT 6.28 38.08 7.48 38.36 ;
  LAYER M2 ;
        RECT 1.12 43.12 2.32 43.4 ;
  LAYER M2 ;
        RECT 2.84 43.12 4.04 43.4 ;
  LAYER M2 ;
        RECT 6.28 45.64 7.48 45.92 ;
  LAYER M2 ;
        RECT 2.15 38.08 3.87 38.36 ;
  LAYER M2 ;
        RECT 4.73 38.08 6.45 38.36 ;
  LAYER M2 ;
        RECT 1.99 38.08 2.31 38.36 ;
  LAYER M1 ;
        RECT 2.025 38.22 2.275 43.26 ;
  LAYER M2 ;
        RECT 1.99 43.12 2.31 43.4 ;
  LAYER M2 ;
        RECT 2.15 43.12 3.01 43.4 ;
  LAYER M2 ;
        RECT 3.71 43.12 4.03 43.4 ;
  LAYER M3 ;
        RECT 3.73 43.26 4.01 45.78 ;
  LAYER M2 ;
        RECT 3.87 45.64 6.45 45.92 ;
  LAYER M1 ;
        RECT 2.025 38.135 2.275 38.305 ;
  LAYER M2 ;
        RECT 1.98 38.08 2.32 38.36 ;
  LAYER M1 ;
        RECT 2.025 43.175 2.275 43.345 ;
  LAYER M2 ;
        RECT 1.98 43.12 2.32 43.4 ;
  LAYER M1 ;
        RECT 2.025 38.135 2.275 38.305 ;
  LAYER M2 ;
        RECT 1.98 38.08 2.32 38.36 ;
  LAYER M1 ;
        RECT 2.025 43.175 2.275 43.345 ;
  LAYER M2 ;
        RECT 1.98 43.12 2.32 43.4 ;
  LAYER M1 ;
        RECT 2.025 38.135 2.275 38.305 ;
  LAYER M2 ;
        RECT 1.98 38.08 2.32 38.36 ;
  LAYER M1 ;
        RECT 2.025 43.175 2.275 43.345 ;
  LAYER M2 ;
        RECT 1.98 43.12 2.32 43.4 ;
  LAYER M1 ;
        RECT 2.025 38.135 2.275 38.305 ;
  LAYER M2 ;
        RECT 1.98 38.08 2.32 38.36 ;
  LAYER M1 ;
        RECT 2.025 43.175 2.275 43.345 ;
  LAYER M2 ;
        RECT 1.98 43.12 2.32 43.4 ;
  LAYER M1 ;
        RECT 2.025 38.135 2.275 38.305 ;
  LAYER M2 ;
        RECT 1.98 38.08 2.32 38.36 ;
  LAYER M1 ;
        RECT 2.025 43.175 2.275 43.345 ;
  LAYER M2 ;
        RECT 1.98 43.12 2.32 43.4 ;
  LAYER M2 ;
        RECT 3.71 43.12 4.03 43.4 ;
  LAYER M3 ;
        RECT 3.73 43.1 4.01 43.42 ;
  LAYER M2 ;
        RECT 3.71 45.64 4.03 45.92 ;
  LAYER M3 ;
        RECT 3.73 45.62 4.01 45.94 ;
  LAYER M1 ;
        RECT 2.025 38.135 2.275 38.305 ;
  LAYER M2 ;
        RECT 1.98 38.08 2.32 38.36 ;
  LAYER M1 ;
        RECT 2.025 43.175 2.275 43.345 ;
  LAYER M2 ;
        RECT 1.98 43.12 2.32 43.4 ;
  LAYER M2 ;
        RECT 3.71 43.12 4.03 43.4 ;
  LAYER M3 ;
        RECT 3.73 43.1 4.01 43.42 ;
  LAYER M2 ;
        RECT 3.71 45.64 4.03 45.92 ;
  LAYER M3 ;
        RECT 3.73 45.62 4.01 45.94 ;
  LAYER M1 ;
        RECT 8.905 43.175 9.155 46.705 ;
  LAYER M1 ;
        RECT 8.905 46.955 9.155 47.965 ;
  LAYER M1 ;
        RECT 8.905 49.055 9.155 50.065 ;
  LAYER M1 ;
        RECT 8.475 43.175 8.725 46.705 ;
  LAYER M1 ;
        RECT 9.335 43.175 9.585 46.705 ;
  LAYER M2 ;
        RECT 8.43 49.42 9.63 49.7 ;
  LAYER M2 ;
        RECT 8.43 43.54 9.63 43.82 ;
  LAYER M2 ;
        RECT 8 43.12 9.2 43.4 ;
  LAYER M2 ;
        RECT 8 47.32 9.2 47.6 ;
  LAYER M3 ;
        RECT 9.32 43.52 9.6 49.72 ;
  LAYER M1 ;
        RECT 8.905 38.975 9.155 42.505 ;
  LAYER M1 ;
        RECT 8.905 37.715 9.155 38.725 ;
  LAYER M1 ;
        RECT 8.905 35.615 9.155 36.625 ;
  LAYER M1 ;
        RECT 8.475 38.975 8.725 42.505 ;
  LAYER M1 ;
        RECT 9.335 38.975 9.585 42.505 ;
  LAYER M2 ;
        RECT 8.43 35.98 9.63 36.26 ;
  LAYER M2 ;
        RECT 8.43 41.86 9.63 42.14 ;
  LAYER M2 ;
        RECT 8 42.28 9.2 42.56 ;
  LAYER M2 ;
        RECT 8 38.08 9.2 38.36 ;
  LAYER M3 ;
        RECT 9.32 35.96 9.6 42.16 ;
  LAYER M1 ;
        RECT 1.165 43.175 1.415 46.705 ;
  LAYER M1 ;
        RECT 1.165 46.955 1.415 47.965 ;
  LAYER M1 ;
        RECT 1.165 49.055 1.415 50.065 ;
  LAYER M1 ;
        RECT 1.595 43.175 1.845 46.705 ;
  LAYER M1 ;
        RECT 0.735 43.175 0.985 46.705 ;
  LAYER M2 ;
        RECT 0.69 49.42 1.89 49.7 ;
  LAYER M2 ;
        RECT 0.69 43.54 1.89 43.82 ;
  LAYER M2 ;
        RECT 1.12 43.12 2.32 43.4 ;
  LAYER M2 ;
        RECT 1.12 47.32 2.32 47.6 ;
  LAYER M3 ;
        RECT 0.72 43.52 1 49.72 ;
  LAYER M1 ;
        RECT 3.745 38.975 3.995 42.505 ;
  LAYER M1 ;
        RECT 3.745 37.715 3.995 38.725 ;
  LAYER M1 ;
        RECT 3.745 35.615 3.995 36.625 ;
  LAYER M1 ;
        RECT 4.175 38.975 4.425 42.505 ;
  LAYER M1 ;
        RECT 3.315 38.975 3.565 42.505 ;
  LAYER M2 ;
        RECT 3.27 35.98 4.47 36.26 ;
  LAYER M2 ;
        RECT 3.27 41.86 4.47 42.14 ;
  LAYER M2 ;
        RECT 3.7 42.28 4.9 42.56 ;
  LAYER M2 ;
        RECT 3.7 38.08 4.9 38.36 ;
  LAYER M3 ;
        RECT 3.3 35.96 3.58 42.16 ;
  LAYER M1 ;
        RECT 6.325 38.975 6.575 42.505 ;
  LAYER M1 ;
        RECT 6.325 37.715 6.575 38.725 ;
  LAYER M1 ;
        RECT 6.325 35.615 6.575 36.625 ;
  LAYER M1 ;
        RECT 6.755 38.975 7.005 42.505 ;
  LAYER M1 ;
        RECT 5.895 38.975 6.145 42.505 ;
  LAYER M2 ;
        RECT 5.85 35.98 7.05 36.26 ;
  LAYER M2 ;
        RECT 5.85 41.86 7.05 42.14 ;
  LAYER M2 ;
        RECT 6.28 42.28 7.48 42.56 ;
  LAYER M2 ;
        RECT 6.28 38.08 7.48 38.36 ;
  LAYER M3 ;
        RECT 5.88 35.96 6.16 42.16 ;
  LAYER M1 ;
        RECT 3.745 43.175 3.995 46.705 ;
  LAYER M1 ;
        RECT 3.745 46.955 3.995 47.965 ;
  LAYER M1 ;
        RECT 3.745 49.055 3.995 50.065 ;
  LAYER M1 ;
        RECT 3.315 43.175 3.565 46.705 ;
  LAYER M1 ;
        RECT 4.175 43.175 4.425 46.705 ;
  LAYER M2 ;
        RECT 3.27 49.42 4.47 49.7 ;
  LAYER M2 ;
        RECT 3.27 43.54 4.47 43.82 ;
  LAYER M2 ;
        RECT 2.84 43.12 4.04 43.4 ;
  LAYER M2 ;
        RECT 2.84 47.32 4.04 47.6 ;
  LAYER M3 ;
        RECT 4.16 43.52 4.44 49.72 ;
  LAYER M1 ;
        RECT 1.165 38.975 1.415 42.505 ;
  LAYER M1 ;
        RECT 1.165 37.715 1.415 38.725 ;
  LAYER M1 ;
        RECT 1.165 35.615 1.415 36.625 ;
  LAYER M1 ;
        RECT 1.595 38.975 1.845 42.505 ;
  LAYER M1 ;
        RECT 0.735 38.975 0.985 42.505 ;
  LAYER M2 ;
        RECT 0.69 35.98 1.89 36.26 ;
  LAYER M2 ;
        RECT 0.69 41.86 1.89 42.14 ;
  LAYER M2 ;
        RECT 1.12 42.28 2.32 42.56 ;
  LAYER M2 ;
        RECT 1.12 38.08 2.32 38.36 ;
  LAYER M3 ;
        RECT 0.72 35.96 1 42.16 ;
  LAYER M1 ;
        RECT 6.325 46.535 6.575 50.065 ;
  LAYER M1 ;
        RECT 6.325 45.275 6.575 46.285 ;
  LAYER M1 ;
        RECT 6.325 43.175 6.575 44.185 ;
  LAYER M1 ;
        RECT 6.755 46.535 7.005 50.065 ;
  LAYER M1 ;
        RECT 5.895 46.535 6.145 50.065 ;
  LAYER M2 ;
        RECT 5.85 43.54 7.05 43.82 ;
  LAYER M2 ;
        RECT 5.85 49.42 7.05 49.7 ;
  LAYER M2 ;
        RECT 6.28 49.84 7.48 50.12 ;
  LAYER M2 ;
        RECT 6.28 45.64 7.48 45.92 ;
  LAYER M3 ;
        RECT 5.88 43.52 6.16 49.72 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 8 17.08 9.2 17.36 ;
  LAYER M2 ;
        RECT 8.01 7.84 8.33 8.12 ;
  LAYER M1 ;
        RECT 8.045 7.98 8.295 17.22 ;
  LAYER M2 ;
        RECT 8.01 17.08 8.33 17.36 ;
  LAYER M2 ;
        RECT 2.15 12.04 3.87 12.32 ;
  LAYER M2 ;
        RECT 4.73 12.04 5.59 12.32 ;
  LAYER M1 ;
        RECT 5.465 12.18 5.715 12.6 ;
  LAYER M2 ;
        RECT 5.59 12.46 8.17 12.74 ;
  LAYER M1 ;
        RECT 8.045 12.515 8.295 12.685 ;
  LAYER M1 ;
        RECT 5.465 12.095 5.715 12.265 ;
  LAYER M2 ;
        RECT 5.42 12.04 5.76 12.32 ;
  LAYER M1 ;
        RECT 5.465 12.515 5.715 12.685 ;
  LAYER M2 ;
        RECT 5.42 12.46 5.76 12.74 ;
  LAYER M1 ;
        RECT 8.045 12.515 8.295 12.685 ;
  LAYER M2 ;
        RECT 8 12.46 8.34 12.74 ;
  LAYER M1 ;
        RECT 5.465 12.095 5.715 12.265 ;
  LAYER M2 ;
        RECT 5.42 12.04 5.76 12.32 ;
  LAYER M1 ;
        RECT 5.465 12.515 5.715 12.685 ;
  LAYER M2 ;
        RECT 5.42 12.46 5.76 12.74 ;
  LAYER M1 ;
        RECT 8.045 12.515 8.295 12.685 ;
  LAYER M2 ;
        RECT 8 12.46 8.34 12.74 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.88 2.32 13.16 ;
  LAYER M2 ;
        RECT 2.84 12.88 4.04 13.16 ;
  LAYER M2 ;
        RECT 6.28 15.4 7.48 15.68 ;
  LAYER M2 ;
        RECT 2.15 7.84 3.87 8.12 ;
  LAYER M2 ;
        RECT 4.73 7.84 6.45 8.12 ;
  LAYER M2 ;
        RECT 1.99 7.84 2.31 8.12 ;
  LAYER M1 ;
        RECT 2.025 7.98 2.275 13.02 ;
  LAYER M2 ;
        RECT 1.99 12.88 2.31 13.16 ;
  LAYER M2 ;
        RECT 2.15 12.88 3.01 13.16 ;
  LAYER M2 ;
        RECT 3.71 12.88 4.03 13.16 ;
  LAYER M3 ;
        RECT 3.73 13.02 4.01 15.54 ;
  LAYER M2 ;
        RECT 3.87 15.4 6.45 15.68 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 12.935 2.275 13.105 ;
  LAYER M2 ;
        RECT 1.98 12.88 2.32 13.16 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 12.935 2.275 13.105 ;
  LAYER M2 ;
        RECT 1.98 12.88 2.32 13.16 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 12.935 2.275 13.105 ;
  LAYER M2 ;
        RECT 1.98 12.88 2.32 13.16 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 12.935 2.275 13.105 ;
  LAYER M2 ;
        RECT 1.98 12.88 2.32 13.16 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 12.935 2.275 13.105 ;
  LAYER M2 ;
        RECT 1.98 12.88 2.32 13.16 ;
  LAYER M2 ;
        RECT 3.71 12.88 4.03 13.16 ;
  LAYER M3 ;
        RECT 3.73 12.86 4.01 13.18 ;
  LAYER M2 ;
        RECT 3.71 15.4 4.03 15.68 ;
  LAYER M3 ;
        RECT 3.73 15.38 4.01 15.7 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.065 ;
  LAYER M2 ;
        RECT 1.98 7.84 2.32 8.12 ;
  LAYER M1 ;
        RECT 2.025 12.935 2.275 13.105 ;
  LAYER M2 ;
        RECT 1.98 12.88 2.32 13.16 ;
  LAYER M2 ;
        RECT 3.71 12.88 4.03 13.16 ;
  LAYER M3 ;
        RECT 3.73 12.86 4.01 13.18 ;
  LAYER M2 ;
        RECT 3.71 15.4 4.03 15.68 ;
  LAYER M3 ;
        RECT 3.73 15.38 4.01 15.7 ;
  LAYER M1 ;
        RECT 8.905 12.935 9.155 16.465 ;
  LAYER M1 ;
        RECT 8.905 16.715 9.155 17.725 ;
  LAYER M1 ;
        RECT 8.905 18.815 9.155 19.825 ;
  LAYER M1 ;
        RECT 8.475 12.935 8.725 16.465 ;
  LAYER M1 ;
        RECT 9.335 12.935 9.585 16.465 ;
  LAYER M2 ;
        RECT 8.43 19.18 9.63 19.46 ;
  LAYER M2 ;
        RECT 8.43 13.3 9.63 13.58 ;
  LAYER M2 ;
        RECT 8 12.88 9.2 13.16 ;
  LAYER M2 ;
        RECT 8 17.08 9.2 17.36 ;
  LAYER M3 ;
        RECT 9.32 13.28 9.6 19.48 ;
  LAYER M1 ;
        RECT 8.905 8.735 9.155 12.265 ;
  LAYER M1 ;
        RECT 8.905 7.475 9.155 8.485 ;
  LAYER M1 ;
        RECT 8.905 5.375 9.155 6.385 ;
  LAYER M1 ;
        RECT 8.475 8.735 8.725 12.265 ;
  LAYER M1 ;
        RECT 9.335 8.735 9.585 12.265 ;
  LAYER M2 ;
        RECT 8.43 5.74 9.63 6.02 ;
  LAYER M2 ;
        RECT 8.43 11.62 9.63 11.9 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M3 ;
        RECT 9.32 5.72 9.6 11.92 ;
  LAYER M1 ;
        RECT 1.165 12.935 1.415 16.465 ;
  LAYER M1 ;
        RECT 1.165 16.715 1.415 17.725 ;
  LAYER M1 ;
        RECT 1.165 18.815 1.415 19.825 ;
  LAYER M1 ;
        RECT 1.595 12.935 1.845 16.465 ;
  LAYER M1 ;
        RECT 0.735 12.935 0.985 16.465 ;
  LAYER M2 ;
        RECT 0.69 19.18 1.89 19.46 ;
  LAYER M2 ;
        RECT 0.69 13.3 1.89 13.58 ;
  LAYER M2 ;
        RECT 1.12 12.88 2.32 13.16 ;
  LAYER M2 ;
        RECT 1.12 17.08 2.32 17.36 ;
  LAYER M3 ;
        RECT 0.72 13.28 1 19.48 ;
  LAYER M1 ;
        RECT 3.745 8.735 3.995 12.265 ;
  LAYER M1 ;
        RECT 3.745 7.475 3.995 8.485 ;
  LAYER M1 ;
        RECT 3.745 5.375 3.995 6.385 ;
  LAYER M1 ;
        RECT 4.175 8.735 4.425 12.265 ;
  LAYER M1 ;
        RECT 3.315 8.735 3.565 12.265 ;
  LAYER M2 ;
        RECT 3.27 5.74 4.47 6.02 ;
  LAYER M2 ;
        RECT 3.27 11.62 4.47 11.9 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M3 ;
        RECT 3.3 5.72 3.58 11.92 ;
  LAYER M1 ;
        RECT 6.325 8.735 6.575 12.265 ;
  LAYER M1 ;
        RECT 6.325 7.475 6.575 8.485 ;
  LAYER M1 ;
        RECT 6.325 5.375 6.575 6.385 ;
  LAYER M1 ;
        RECT 6.755 8.735 7.005 12.265 ;
  LAYER M1 ;
        RECT 5.895 8.735 6.145 12.265 ;
  LAYER M2 ;
        RECT 5.85 5.74 7.05 6.02 ;
  LAYER M2 ;
        RECT 5.85 11.62 7.05 11.9 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M3 ;
        RECT 5.88 5.72 6.16 11.92 ;
  LAYER M1 ;
        RECT 3.745 12.935 3.995 16.465 ;
  LAYER M1 ;
        RECT 3.745 16.715 3.995 17.725 ;
  LAYER M1 ;
        RECT 3.745 18.815 3.995 19.825 ;
  LAYER M1 ;
        RECT 3.315 12.935 3.565 16.465 ;
  LAYER M1 ;
        RECT 4.175 12.935 4.425 16.465 ;
  LAYER M2 ;
        RECT 3.27 19.18 4.47 19.46 ;
  LAYER M2 ;
        RECT 3.27 13.3 4.47 13.58 ;
  LAYER M2 ;
        RECT 2.84 12.88 4.04 13.16 ;
  LAYER M2 ;
        RECT 2.84 17.08 4.04 17.36 ;
  LAYER M3 ;
        RECT 4.16 13.28 4.44 19.48 ;
  LAYER M1 ;
        RECT 1.165 8.735 1.415 12.265 ;
  LAYER M1 ;
        RECT 1.165 7.475 1.415 8.485 ;
  LAYER M1 ;
        RECT 1.165 5.375 1.415 6.385 ;
  LAYER M1 ;
        RECT 1.595 8.735 1.845 12.265 ;
  LAYER M1 ;
        RECT 0.735 8.735 0.985 12.265 ;
  LAYER M2 ;
        RECT 0.69 5.74 1.89 6.02 ;
  LAYER M2 ;
        RECT 0.69 11.62 1.89 11.9 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M3 ;
        RECT 0.72 5.72 1 11.92 ;
  LAYER M1 ;
        RECT 6.325 16.295 6.575 19.825 ;
  LAYER M1 ;
        RECT 6.325 15.035 6.575 16.045 ;
  LAYER M1 ;
        RECT 6.325 12.935 6.575 13.945 ;
  LAYER M1 ;
        RECT 6.755 16.295 7.005 19.825 ;
  LAYER M1 ;
        RECT 5.895 16.295 6.145 19.825 ;
  LAYER M2 ;
        RECT 5.85 13.3 7.05 13.58 ;
  LAYER M2 ;
        RECT 5.85 19.18 7.05 19.46 ;
  LAYER M2 ;
        RECT 6.28 19.6 7.48 19.88 ;
  LAYER M2 ;
        RECT 6.28 15.4 7.48 15.68 ;
  LAYER M3 ;
        RECT 5.88 13.28 6.16 19.48 ;
  LAYER M2 ;
        RECT 1.12 27.16 2.32 27.44 ;
  LAYER M2 ;
        RECT 3.7 27.16 4.9 27.44 ;
  LAYER M2 ;
        RECT 8 22.96 9.2 23.24 ;
  LAYER M2 ;
        RECT 8 32.2 9.2 32.48 ;
  LAYER M2 ;
        RECT 8.01 22.96 8.33 23.24 ;
  LAYER M1 ;
        RECT 8.045 23.1 8.295 32.34 ;
  LAYER M2 ;
        RECT 8.01 32.2 8.33 32.48 ;
  LAYER M2 ;
        RECT 2.15 27.16 3.87 27.44 ;
  LAYER M2 ;
        RECT 4.73 27.16 5.59 27.44 ;
  LAYER M1 ;
        RECT 5.465 27.3 5.715 27.72 ;
  LAYER M2 ;
        RECT 5.59 27.58 8.17 27.86 ;
  LAYER M1 ;
        RECT 8.045 27.635 8.295 27.805 ;
  LAYER M1 ;
        RECT 5.465 27.215 5.715 27.385 ;
  LAYER M2 ;
        RECT 5.42 27.16 5.76 27.44 ;
  LAYER M1 ;
        RECT 5.465 27.635 5.715 27.805 ;
  LAYER M2 ;
        RECT 5.42 27.58 5.76 27.86 ;
  LAYER M1 ;
        RECT 8.045 27.635 8.295 27.805 ;
  LAYER M2 ;
        RECT 8 27.58 8.34 27.86 ;
  LAYER M1 ;
        RECT 5.465 27.215 5.715 27.385 ;
  LAYER M2 ;
        RECT 5.42 27.16 5.76 27.44 ;
  LAYER M1 ;
        RECT 5.465 27.635 5.715 27.805 ;
  LAYER M2 ;
        RECT 5.42 27.58 5.76 27.86 ;
  LAYER M1 ;
        RECT 8.045 27.635 8.295 27.805 ;
  LAYER M2 ;
        RECT 8 27.58 8.34 27.86 ;
  LAYER M2 ;
        RECT 1.12 22.96 2.32 23.24 ;
  LAYER M2 ;
        RECT 3.7 22.96 4.9 23.24 ;
  LAYER M2 ;
        RECT 6.28 22.96 7.48 23.24 ;
  LAYER M2 ;
        RECT 1.12 28 2.32 28.28 ;
  LAYER M2 ;
        RECT 2.84 28 4.04 28.28 ;
  LAYER M2 ;
        RECT 6.28 30.52 7.48 30.8 ;
  LAYER M2 ;
        RECT 2.15 22.96 3.87 23.24 ;
  LAYER M2 ;
        RECT 4.73 22.96 6.45 23.24 ;
  LAYER M2 ;
        RECT 1.99 22.96 2.31 23.24 ;
  LAYER M1 ;
        RECT 2.025 23.1 2.275 28.14 ;
  LAYER M2 ;
        RECT 1.99 28 2.31 28.28 ;
  LAYER M2 ;
        RECT 2.15 28 3.01 28.28 ;
  LAYER M2 ;
        RECT 3.71 28 4.03 28.28 ;
  LAYER M3 ;
        RECT 3.73 28.14 4.01 30.66 ;
  LAYER M2 ;
        RECT 3.87 30.52 6.45 30.8 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 23.185 ;
  LAYER M2 ;
        RECT 1.98 22.96 2.32 23.24 ;
  LAYER M1 ;
        RECT 2.025 28.055 2.275 28.225 ;
  LAYER M2 ;
        RECT 1.98 28 2.32 28.28 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 23.185 ;
  LAYER M2 ;
        RECT 1.98 22.96 2.32 23.24 ;
  LAYER M1 ;
        RECT 2.025 28.055 2.275 28.225 ;
  LAYER M2 ;
        RECT 1.98 28 2.32 28.28 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 23.185 ;
  LAYER M2 ;
        RECT 1.98 22.96 2.32 23.24 ;
  LAYER M1 ;
        RECT 2.025 28.055 2.275 28.225 ;
  LAYER M2 ;
        RECT 1.98 28 2.32 28.28 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 23.185 ;
  LAYER M2 ;
        RECT 1.98 22.96 2.32 23.24 ;
  LAYER M1 ;
        RECT 2.025 28.055 2.275 28.225 ;
  LAYER M2 ;
        RECT 1.98 28 2.32 28.28 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 23.185 ;
  LAYER M2 ;
        RECT 1.98 22.96 2.32 23.24 ;
  LAYER M1 ;
        RECT 2.025 28.055 2.275 28.225 ;
  LAYER M2 ;
        RECT 1.98 28 2.32 28.28 ;
  LAYER M2 ;
        RECT 3.71 28 4.03 28.28 ;
  LAYER M3 ;
        RECT 3.73 27.98 4.01 28.3 ;
  LAYER M2 ;
        RECT 3.71 30.52 4.03 30.8 ;
  LAYER M3 ;
        RECT 3.73 30.5 4.01 30.82 ;
  LAYER M1 ;
        RECT 2.025 23.015 2.275 23.185 ;
  LAYER M2 ;
        RECT 1.98 22.96 2.32 23.24 ;
  LAYER M1 ;
        RECT 2.025 28.055 2.275 28.225 ;
  LAYER M2 ;
        RECT 1.98 28 2.32 28.28 ;
  LAYER M2 ;
        RECT 3.71 28 4.03 28.28 ;
  LAYER M3 ;
        RECT 3.73 27.98 4.01 28.3 ;
  LAYER M2 ;
        RECT 3.71 30.52 4.03 30.8 ;
  LAYER M3 ;
        RECT 3.73 30.5 4.01 30.82 ;
  LAYER M1 ;
        RECT 8.905 28.055 9.155 31.585 ;
  LAYER M1 ;
        RECT 8.905 31.835 9.155 32.845 ;
  LAYER M1 ;
        RECT 8.905 33.935 9.155 34.945 ;
  LAYER M1 ;
        RECT 8.475 28.055 8.725 31.585 ;
  LAYER M1 ;
        RECT 9.335 28.055 9.585 31.585 ;
  LAYER M2 ;
        RECT 8.43 34.3 9.63 34.58 ;
  LAYER M2 ;
        RECT 8.43 28.42 9.63 28.7 ;
  LAYER M2 ;
        RECT 8 28 9.2 28.28 ;
  LAYER M2 ;
        RECT 8 32.2 9.2 32.48 ;
  LAYER M3 ;
        RECT 9.32 28.4 9.6 34.6 ;
  LAYER M1 ;
        RECT 8.905 23.855 9.155 27.385 ;
  LAYER M1 ;
        RECT 8.905 22.595 9.155 23.605 ;
  LAYER M1 ;
        RECT 8.905 20.495 9.155 21.505 ;
  LAYER M1 ;
        RECT 8.475 23.855 8.725 27.385 ;
  LAYER M1 ;
        RECT 9.335 23.855 9.585 27.385 ;
  LAYER M2 ;
        RECT 8.43 20.86 9.63 21.14 ;
  LAYER M2 ;
        RECT 8.43 26.74 9.63 27.02 ;
  LAYER M2 ;
        RECT 8 27.16 9.2 27.44 ;
  LAYER M2 ;
        RECT 8 22.96 9.2 23.24 ;
  LAYER M3 ;
        RECT 9.32 20.84 9.6 27.04 ;
  LAYER M1 ;
        RECT 1.165 28.055 1.415 31.585 ;
  LAYER M1 ;
        RECT 1.165 31.835 1.415 32.845 ;
  LAYER M1 ;
        RECT 1.165 33.935 1.415 34.945 ;
  LAYER M1 ;
        RECT 1.595 28.055 1.845 31.585 ;
  LAYER M1 ;
        RECT 0.735 28.055 0.985 31.585 ;
  LAYER M2 ;
        RECT 0.69 34.3 1.89 34.58 ;
  LAYER M2 ;
        RECT 0.69 28.42 1.89 28.7 ;
  LAYER M2 ;
        RECT 1.12 28 2.32 28.28 ;
  LAYER M2 ;
        RECT 1.12 32.2 2.32 32.48 ;
  LAYER M3 ;
        RECT 0.72 28.4 1 34.6 ;
  LAYER M1 ;
        RECT 3.745 23.855 3.995 27.385 ;
  LAYER M1 ;
        RECT 3.745 22.595 3.995 23.605 ;
  LAYER M1 ;
        RECT 3.745 20.495 3.995 21.505 ;
  LAYER M1 ;
        RECT 4.175 23.855 4.425 27.385 ;
  LAYER M1 ;
        RECT 3.315 23.855 3.565 27.385 ;
  LAYER M2 ;
        RECT 3.27 20.86 4.47 21.14 ;
  LAYER M2 ;
        RECT 3.27 26.74 4.47 27.02 ;
  LAYER M2 ;
        RECT 3.7 27.16 4.9 27.44 ;
  LAYER M2 ;
        RECT 3.7 22.96 4.9 23.24 ;
  LAYER M3 ;
        RECT 3.3 20.84 3.58 27.04 ;
  LAYER M1 ;
        RECT 6.325 23.855 6.575 27.385 ;
  LAYER M1 ;
        RECT 6.325 22.595 6.575 23.605 ;
  LAYER M1 ;
        RECT 6.325 20.495 6.575 21.505 ;
  LAYER M1 ;
        RECT 6.755 23.855 7.005 27.385 ;
  LAYER M1 ;
        RECT 5.895 23.855 6.145 27.385 ;
  LAYER M2 ;
        RECT 5.85 20.86 7.05 21.14 ;
  LAYER M2 ;
        RECT 5.85 26.74 7.05 27.02 ;
  LAYER M2 ;
        RECT 6.28 27.16 7.48 27.44 ;
  LAYER M2 ;
        RECT 6.28 22.96 7.48 23.24 ;
  LAYER M3 ;
        RECT 5.88 20.84 6.16 27.04 ;
  LAYER M1 ;
        RECT 3.745 28.055 3.995 31.585 ;
  LAYER M1 ;
        RECT 3.745 31.835 3.995 32.845 ;
  LAYER M1 ;
        RECT 3.745 33.935 3.995 34.945 ;
  LAYER M1 ;
        RECT 3.315 28.055 3.565 31.585 ;
  LAYER M1 ;
        RECT 4.175 28.055 4.425 31.585 ;
  LAYER M2 ;
        RECT 3.27 34.3 4.47 34.58 ;
  LAYER M2 ;
        RECT 3.27 28.42 4.47 28.7 ;
  LAYER M2 ;
        RECT 2.84 28 4.04 28.28 ;
  LAYER M2 ;
        RECT 2.84 32.2 4.04 32.48 ;
  LAYER M3 ;
        RECT 4.16 28.4 4.44 34.6 ;
  LAYER M1 ;
        RECT 1.165 23.855 1.415 27.385 ;
  LAYER M1 ;
        RECT 1.165 22.595 1.415 23.605 ;
  LAYER M1 ;
        RECT 1.165 20.495 1.415 21.505 ;
  LAYER M1 ;
        RECT 1.595 23.855 1.845 27.385 ;
  LAYER M1 ;
        RECT 0.735 23.855 0.985 27.385 ;
  LAYER M2 ;
        RECT 0.69 20.86 1.89 21.14 ;
  LAYER M2 ;
        RECT 0.69 26.74 1.89 27.02 ;
  LAYER M2 ;
        RECT 1.12 27.16 2.32 27.44 ;
  LAYER M2 ;
        RECT 1.12 22.96 2.32 23.24 ;
  LAYER M3 ;
        RECT 0.72 20.84 1 27.04 ;
  LAYER M1 ;
        RECT 6.325 31.415 6.575 34.945 ;
  LAYER M1 ;
        RECT 6.325 30.155 6.575 31.165 ;
  LAYER M1 ;
        RECT 6.325 28.055 6.575 29.065 ;
  LAYER M1 ;
        RECT 6.755 31.415 7.005 34.945 ;
  LAYER M1 ;
        RECT 5.895 31.415 6.145 34.945 ;
  LAYER M2 ;
        RECT 5.85 28.42 7.05 28.7 ;
  LAYER M2 ;
        RECT 5.85 34.3 7.05 34.58 ;
  LAYER M2 ;
        RECT 6.28 34.72 7.48 35 ;
  LAYER M2 ;
        RECT 6.28 30.52 7.48 30.8 ;
  LAYER M3 ;
        RECT 5.88 28.4 6.16 34.6 ;
  LAYER M4 ;
        RECT 11.18 1.93 19.48 10.23 ;
  LAYER M4 ;
        RECT 19.03 1.46 19.48 3.98 ;
  LAYER M5 ;
        RECT 11.405 9.25 11.855 11.77 ;
  LAYER M4 ;
        RECT 10.585 10.94 19.515 11.74 ;
  LAYER M4 ;
        RECT 10.585 0.86 19.515 1.66 ;
  LAYER M4 ;
        RECT 11.18 14.53 19.48 22.83 ;
  LAYER M4 ;
        RECT 19.03 14.06 19.48 16.58 ;
  LAYER M5 ;
        RECT 11.405 21.85 11.855 24.37 ;
  LAYER M4 ;
        RECT 10.585 23.54 19.515 24.34 ;
  LAYER M4 ;
        RECT 10.585 13.46 19.515 14.26 ;
  LAYER M4 ;
        RECT 11.18 27.13 19.48 35.43 ;
  LAYER M4 ;
        RECT 19.03 26.66 19.48 29.18 ;
  LAYER M5 ;
        RECT 11.405 34.45 11.855 36.97 ;
  LAYER M4 ;
        RECT 10.585 36.14 19.515 36.94 ;
  LAYER M4 ;
        RECT 10.585 26.06 19.515 26.86 ;
  LAYER M4 ;
        RECT 11.18 39.73 19.48 48.03 ;
  LAYER M4 ;
        RECT 19.03 39.26 19.48 41.78 ;
  LAYER M5 ;
        RECT 11.405 47.05 11.855 49.57 ;
  LAYER M4 ;
        RECT 10.585 48.74 19.515 49.54 ;
  LAYER M4 ;
        RECT 10.585 38.66 19.515 39.46 ;
  END 
END TWO_BIT_RES_DAC
